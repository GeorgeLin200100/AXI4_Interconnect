`ifndef TOP_DEFINES_SVH
`define TOP_DEFINES_SVH

    `define SLAVE_ADDR_REGION_SIZE  32'h00FF_FFFF
    `define SLAVE_0_BASE_ADDR       32'h0000_0000
    `define SLAVE_1_BASE_ADDR       32'h0100_0000
    `define SLAVE_2_BASE_ADDR       32'h0200_0000
    `define SLAVE_3_BASE_ADDR       32'h0300_0000

`endif