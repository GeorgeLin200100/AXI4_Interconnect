//
`resetall
`timescale 1ns / 1ps
`default_nettype none
`include "axi_tmr_signal_define.vh"

module axi_tmr_voter_ds #
(
    // Width of data bus in bits
    parameter DATA_WIDTH = 64,
    // Width of address bus in bits
    parameter ADDR_WIDTH = 32,
    // Width of wstrb (width of data bus in words)
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    // Input ID field width (from AXI masters)
    parameter S_ID_WIDTH = 8,
    // Output ID field width (towards AXI slaves)
    // Additional bits required for response routing
    parameter M_ID_WIDTH = S_ID_WIDTH+$clog2(3),
    // Propagate awuser signal
    parameter AWUSER_ENABLE = 0,
    // Width of awuser signal
    parameter AWUSER_WIDTH = 1,
    // Propagate wuser signal
    parameter WUSER_ENABLE = 0,
    // Width of wuser signal
    parameter WUSER_WIDTH = 1,
    // Propagate buser signal
    parameter BUSER_ENABLE = 0,
    // Width of buser signal
    parameter BUSER_WIDTH = 1,
    // Propagate aruser signal
    parameter ARUSER_ENABLE = 0,
    // Width of aruser signal
    parameter ARUSER_WIDTH = 1,
    // Propagate ruser signal
    parameter RUSER_ENABLE = 0,
    // Width of ruser signal
    parameter RUSER_WIDTH = 1,
    // Number of concurrent unique IDs
    parameter S00_THREADS = 8,
    // Number of concurrent operations
    parameter S00_ACCEPT = 16,
    // Number of concurrent unique IDs
    parameter S01_THREADS = 8,
    // Number of concurrent operations
    parameter S01_ACCEPT = 16,
    // Number of concurrent unique IDs
    parameter S02_THREADS = 8,
    // Number of concurrent operations
    parameter S02_ACCEPT = 16,
    // Number of regions per master interface
    parameter M_REGIONS = 1,
    // Master interface base addresses
    // M_REGIONS concatenated fields of ADDR_WIDTH bits
    parameter M00_BASE_ADDR = 0, // enable default mapping
    // Master interface address widths
    // M_REGIONS concatenated fields of 32 bits
    parameter M00_ADDR_WIDTH = {M_REGIONS{32'd24}},
    // Read connections between interfaces
    // S_COUNT bits
    parameter M00_CONNECT_READ = 3'b100,  // Slave 0 only connect to Master 2
    // Write connections between interfaces
    // S_COUNT bits
    parameter M00_CONNECT_WRITE = 3'b100, // Slave 0 only connect to Master 2
    // Number of concurrent operations for each master interface
    parameter M00_ISSUE = 8,
    // Secure master (fail operations based on awprot/arprot)
    parameter M00_SECURE = 1, //Slave 0 is secure
    // Master interface base addresses
    // M_REGIONS concatenated fields of ADDR_WIDTH bits
    parameter M01_BASE_ADDR = 0, // enable default mapping
    // Master interface address widths
    // M_REGIONS concatenated fields of 32 bits
    parameter M01_ADDR_WIDTH = {M_REGIONS{32'd24}},
    // Read connections between interfaces
    // S_COUNT bits
    parameter M01_CONNECT_READ = 3'b011, // Slave 1 only connect to Master 0,1
    // Write connections between interfaces
    // S_COUNT bits
    parameter M01_CONNECT_WRITE = 3'b011, // Slave 1 only connect to Master 0,1
    // Number of concurrent operations for each master interface
    parameter M01_ISSUE = 8,
    // Secure master (fail operations based on awprot/arprot)
    parameter M01_SECURE = 0, // Slave 1 is unsecure
    // Master interface base addresses
    // M_REGIONS concatenated fields of ADDR_WIDTH bits
    parameter M02_BASE_ADDR = 0, // enable default mapping
    // Master interface address widths
    // M_REGIONS concatenated fields of 32 bits
    parameter M02_ADDR_WIDTH = {M_REGIONS{32'd24}},
    // Read connections between interfaces
    // S_COUNT bits
    parameter M02_CONNECT_READ = 3'b100, // Slave 2 only connect to Master 2
    // Write connections between interfaces
    // S_COUNT bits
    parameter M02_CONNECT_WRITE = 3'b100, // Slave 2 only connect to Master 2
    // Number of concurrent operations for each master interface
    parameter M02_ISSUE = 8,
    // Secure master (fail operations based on awprot/arprot)
    parameter M02_SECURE = 1,
    // Master interface base addresses
    // M_REGIONS concatenated fields of ADDR_WIDTH bits
    parameter M03_BASE_ADDR = 0,
    // Master interface address widths
    // M_REGIONS concatenated fields of 32 bits
    parameter M03_ADDR_WIDTH = {M_REGIONS{32'd24}},
    // Read connections between interfaces
    // S_COUNT bits
    parameter M03_CONNECT_READ = 3'b011,
    // Write connections between interfaces
    // S_COUNT bits
    parameter M03_CONNECT_WRITE = 3'b011,
    // Number of concurrent operations for each master interface
    parameter M03_ISSUE = 8,
    // Secure master (fail operations based on awprot/arprot)
    parameter M03_SECURE = 0,
    // Slave interface AW channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S00_AW_REG_TYPE = 0,
    // Slave interface W channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S00_W_REG_TYPE = 0,
    // Slave interface B channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S00_B_REG_TYPE = 1,
    // Slave interface AR channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S00_AR_REG_TYPE = 0,
    // Slave interface R channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S00_R_REG_TYPE = 2,
    // Slave interface AW channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S01_AW_REG_TYPE = 0,
    // Slave interface W channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S01_W_REG_TYPE = 0,
    // Slave interface B channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S01_B_REG_TYPE = 1,
    // Slave interface AR channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S01_AR_REG_TYPE = 0,
    // Slave interface R channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S01_R_REG_TYPE = 2,
    // Slave interface AW channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S02_AW_REG_TYPE = 0,
    // Slave interface W channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S02_W_REG_TYPE = 0,
    // Slave interface B channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S02_B_REG_TYPE = 1,
    // Slave interface AR channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S02_AR_REG_TYPE = 0,
    // Slave interface R channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter S02_R_REG_TYPE = 2,
    // Master interface AW channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M00_AW_REG_TYPE = 1,
    // Master interface W channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M00_W_REG_TYPE = 2,
    // Master interface B channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M00_B_REG_TYPE = 0,
    // Master interface AR channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M00_AR_REG_TYPE = 1,
    // Master interface R channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M00_R_REG_TYPE = 0,
    // Master interface AW channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M01_AW_REG_TYPE = 1,
    // Master interface W channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M01_W_REG_TYPE = 2,
    // Master interface B channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M01_B_REG_TYPE = 0,
    // Master interface AR channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M01_AR_REG_TYPE = 1,
    // Master interface R channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M01_R_REG_TYPE = 0,
    // Master interface AW channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M02_AW_REG_TYPE = 1,
    // Master interface W channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M02_W_REG_TYPE = 2,
    // Master interface B channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M02_B_REG_TYPE = 0,
    // Master interface AR channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M02_AR_REG_TYPE = 1,
    // Master interface R channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M02_R_REG_TYPE = 0,
    // Master interface AW channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M03_AW_REG_TYPE = 1,
    // Master interface W channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M03_W_REG_TYPE = 2,
    // Master interface B channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M03_B_REG_TYPE = 0,
    // Master interface AR channel register type (output)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M03_AR_REG_TYPE = 1,
    // Master interface R channel register type (input)
    // 0 to bypass, 1 for simple buffer, 2 for skid buffer
    parameter M03_R_REG_TYPE = 0
)
(
    input  wire                     clk,
    input  wire                     rst,

/* AXI slave interface 
*/
//vd0
    output wire [M_ID_WIDTH-1:0]    s00_vd0_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s00_vd0_axi_awaddr,
    output wire [7:0]               s00_vd0_axi_awlen,
    output wire [2:0]               s00_vd0_axi_awsize,
    output wire [1:0]               s00_vd0_axi_awburst,
    output wire                     s00_vd0_axi_awlock,
    output wire [3:0]               s00_vd0_axi_awcache,
    output wire [2:0]               s00_vd0_axi_awprot,
    output wire [3:0]               s00_vd0_axi_awqos,
    output wire [3:0]               s00_vd0_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s00_vd0_axi_awuser,
    output wire                     s00_vd0_axi_awvalid,
    input  wire                     s00_vd0_axi_awready,
    output wire [DATA_WIDTH-1:0]    s00_vd0_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s00_vd0_axi_wstrb,
    output wire                     s00_vd0_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s00_vd0_axi_wuser,
    output wire                     s00_vd0_axi_wvalid,
    input  wire                     s00_vd0_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd0_axi_bid,
    input  wire [1:0]               s00_vd0_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s00_vd0_axi_buser,
    input  wire                     s00_vd0_axi_bvalid,
    output wire                     s00_vd0_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s00_vd0_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s00_vd0_axi_araddr,
    output wire [7:0]               s00_vd0_axi_arlen,
    output wire [2:0]               s00_vd0_axi_arsize,
    output wire [1:0]               s00_vd0_axi_arburst,
    output wire                     s00_vd0_axi_arlock,
    output wire [3:0]               s00_vd0_axi_arcache,
    output wire [2:0]               s00_vd0_axi_arprot,
    output wire [3:0]               s00_vd0_axi_arqos,
    output wire [3:0]               s00_vd0_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s00_vd0_axi_aruser,
    output wire                     s00_vd0_axi_arvalid,
    input  wire                     s00_vd0_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd0_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s00_vd0_axi_rdata,
    input  wire [1:0]               s00_vd0_axi_rresp,
    input  wire                     s00_vd0_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s00_vd0_axi_ruser,
    input  wire                     s00_vd0_axi_rvalid,
    output wire                     s00_vd0_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s01_vd0_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s01_vd0_axi_awaddr,
    output wire [7:0]               s01_vd0_axi_awlen,
    output wire [2:0]               s01_vd0_axi_awsize,
    output wire [1:0]               s01_vd0_axi_awburst,
    output wire                     s01_vd0_axi_awlock,
    output wire [3:0]               s01_vd0_axi_awcache,
    output wire [2:0]               s01_vd0_axi_awprot,
    output wire [3:0]               s01_vd0_axi_awqos,
    output wire [3:0]               s01_vd0_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s01_vd0_axi_awuser,
    output wire                     s01_vd0_axi_awvalid,
    input  wire                     s01_vd0_axi_awready,
    output wire [DATA_WIDTH-1:0]    s01_vd0_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s01_vd0_axi_wstrb,
    output wire                     s01_vd0_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s01_vd0_axi_wuser,
    output wire                     s01_vd0_axi_wvalid,
    input  wire                     s01_vd0_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd0_axi_bid,
    input  wire [1:0]               s01_vd0_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s01_vd0_axi_buser,
    input  wire                     s01_vd0_axi_bvalid,
    output wire                     s01_vd0_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s01_vd0_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s01_vd0_axi_araddr,
    output wire [7:0]               s01_vd0_axi_arlen,
    output wire [2:0]               s01_vd0_axi_arsize,
    output wire [1:0]               s01_vd0_axi_arburst,
    output wire                     s01_vd0_axi_arlock,
    output wire [3:0]               s01_vd0_axi_arcache,
    output wire [2:0]               s01_vd0_axi_arprot,
    output wire [3:0]               s01_vd0_axi_arqos,
    output wire [3:0]               s01_vd0_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s01_vd0_axi_aruser,
    output wire                     s01_vd0_axi_arvalid,
    input  wire                     s01_vd0_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd0_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s01_vd0_axi_rdata,
    input  wire [1:0]               s01_vd0_axi_rresp,
    input  wire                     s01_vd0_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s01_vd0_axi_ruser,
    input  wire                     s01_vd0_axi_rvalid,
    output wire                     s01_vd0_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s02_vd0_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s02_vd0_axi_awaddr,
    output wire [7:0]               s02_vd0_axi_awlen,
    output wire [2:0]               s02_vd0_axi_awsize,
    output wire [1:0]               s02_vd0_axi_awburst,
    output wire                     s02_vd0_axi_awlock,
    output wire [3:0]               s02_vd0_axi_awcache,
    output wire [2:0]               s02_vd0_axi_awprot,
    output wire [3:0]               s02_vd0_axi_awqos,
    output wire [3:0]               s02_vd0_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s02_vd0_axi_awuser,
    output wire                     s02_vd0_axi_awvalid,
    input  wire                     s02_vd0_axi_awready,
    output wire [DATA_WIDTH-1:0]    s02_vd0_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s02_vd0_axi_wstrb,
    output wire                     s02_vd0_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s02_vd0_axi_wuser,
    output wire                     s02_vd0_axi_wvalid,
    input  wire                     s02_vd0_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd0_axi_bid,
    input  wire [1:0]               s02_vd0_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s02_vd0_axi_buser,
    input  wire                     s02_vd0_axi_bvalid,
    output wire                     s02_vd0_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s02_vd0_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s02_vd0_axi_araddr,
    output wire [7:0]               s02_vd0_axi_arlen,
    output wire [2:0]               s02_vd0_axi_arsize,
    output wire [1:0]               s02_vd0_axi_arburst,
    output wire                     s02_vd0_axi_arlock,
    output wire [3:0]               s02_vd0_axi_arcache,
    output wire [2:0]               s02_vd0_axi_arprot,
    output wire [3:0]               s02_vd0_axi_arqos,
    output wire [3:0]               s02_vd0_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s02_vd0_axi_aruser,
    output wire                     s02_vd0_axi_arvalid,
    input  wire                     s02_vd0_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd0_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s02_vd0_axi_rdata,
    input  wire [1:0]               s02_vd0_axi_rresp,
    input  wire                     s02_vd0_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s02_vd0_axi_ruser,
    input  wire                     s02_vd0_axi_rvalid,
    output wire                     s02_vd0_axi_rready,
//vd1
    output wire [M_ID_WIDTH-1:0]    s00_vd1_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s00_vd1_axi_awaddr,
    output wire [7:0]               s00_vd1_axi_awlen,
    output wire [2:0]               s00_vd1_axi_awsize,
    output wire [1:0]               s00_vd1_axi_awburst,
    output wire                     s00_vd1_axi_awlock,
    output wire [3:0]               s00_vd1_axi_awcache,
    output wire [2:0]               s00_vd1_axi_awprot,
    output wire [3:0]               s00_vd1_axi_awqos,
    output wire [3:0]               s00_vd1_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s00_vd1_axi_awuser,
    output wire                     s00_vd1_axi_awvalid,
    input  wire                     s00_vd1_axi_awready,
    output wire [DATA_WIDTH-1:0]    s00_vd1_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s00_vd1_axi_wstrb,
    output wire                     s00_vd1_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s00_vd1_axi_wuser,
    output wire                     s00_vd1_axi_wvalid,
    input  wire                     s00_vd1_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd1_axi_bid,
    input  wire [1:0]               s00_vd1_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s00_vd1_axi_buser,
    input  wire                     s00_vd1_axi_bvalid,
    output wire                     s00_vd1_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s00_vd1_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s00_vd1_axi_araddr,
    output wire [7:0]               s00_vd1_axi_arlen,
    output wire [2:0]               s00_vd1_axi_arsize,
    output wire [1:0]               s00_vd1_axi_arburst,
    output wire                     s00_vd1_axi_arlock,
    output wire [3:0]               s00_vd1_axi_arcache,
    output wire [2:0]               s00_vd1_axi_arprot,
    output wire [3:0]               s00_vd1_axi_arqos,
    output wire [3:0]               s00_vd1_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s00_vd1_axi_aruser,
    output wire                     s00_vd1_axi_arvalid,
    input  wire                     s00_vd1_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd1_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s00_vd1_axi_rdata,
    input  wire [1:0]               s00_vd1_axi_rresp,
    input  wire                     s00_vd1_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s00_vd1_axi_ruser,
    input  wire                     s00_vd1_axi_rvalid,
    output wire                     s00_vd1_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s01_vd1_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s01_vd1_axi_awaddr,
    output wire [7:0]               s01_vd1_axi_awlen,
    output wire [2:0]               s01_vd1_axi_awsize,
    output wire [1:0]               s01_vd1_axi_awburst,
    output wire                     s01_vd1_axi_awlock,
    output wire [3:0]               s01_vd1_axi_awcache,
    output wire [2:0]               s01_vd1_axi_awprot,
    output wire [3:0]               s01_vd1_axi_awqos,
    output wire [3:0]               s01_vd1_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s01_vd1_axi_awuser,
    output wire                     s01_vd1_axi_awvalid,
    input  wire                     s01_vd1_axi_awready,
    output wire [DATA_WIDTH-1:0]    s01_vd1_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s01_vd1_axi_wstrb,
    output wire                     s01_vd1_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s01_vd1_axi_wuser,
    output wire                     s01_vd1_axi_wvalid,
    input  wire                     s01_vd1_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd1_axi_bid,
    input  wire [1:0]               s01_vd1_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s01_vd1_axi_buser,
    input  wire                     s01_vd1_axi_bvalid,
    output wire                     s01_vd1_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s01_vd1_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s01_vd1_axi_araddr,
    output wire [7:0]               s01_vd1_axi_arlen,
    output wire [2:0]               s01_vd1_axi_arsize,
    output wire [1:0]               s01_vd1_axi_arburst,
    output wire                     s01_vd1_axi_arlock,
    output wire [3:0]               s01_vd1_axi_arcache,
    output wire [2:0]               s01_vd1_axi_arprot,
    output wire [3:0]               s01_vd1_axi_arqos,
    output wire [3:0]               s01_vd1_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s01_vd1_axi_aruser,
    output wire                     s01_vd1_axi_arvalid,
    input  wire                     s01_vd1_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd1_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s01_vd1_axi_rdata,
    input  wire [1:0]               s01_vd1_axi_rresp,
    input  wire                     s01_vd1_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s01_vd1_axi_ruser,
    input  wire                     s01_vd1_axi_rvalid,
    output wire                     s01_vd1_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s02_vd1_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s02_vd1_axi_awaddr,
    output wire [7:0]               s02_vd1_axi_awlen,
    output wire [2:0]               s02_vd1_axi_awsize,
    output wire [1:0]               s02_vd1_axi_awburst,
    output wire                     s02_vd1_axi_awlock,
    output wire [3:0]               s02_vd1_axi_awcache,
    output wire [2:0]               s02_vd1_axi_awprot,
    output wire [3:0]               s02_vd1_axi_awqos,
    output wire [3:0]               s02_vd1_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s02_vd1_axi_awuser,
    output wire                     s02_vd1_axi_awvalid,
    input  wire                     s02_vd1_axi_awready,
    output wire [DATA_WIDTH-1:0]    s02_vd1_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s02_vd1_axi_wstrb,
    output wire                     s02_vd1_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s02_vd1_axi_wuser,
    output wire                     s02_vd1_axi_wvalid,
    input  wire                     s02_vd1_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd1_axi_bid,
    input  wire [1:0]               s02_vd1_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s02_vd1_axi_buser,
    input  wire                     s02_vd1_axi_bvalid,
    output wire                     s02_vd1_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s02_vd1_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s02_vd1_axi_araddr,
    output wire [7:0]               s02_vd1_axi_arlen,
    output wire [2:0]               s02_vd1_axi_arsize,
    output wire [1:0]               s02_vd1_axi_arburst,
    output wire                     s02_vd1_axi_arlock,
    output wire [3:0]               s02_vd1_axi_arcache,
    output wire [2:0]               s02_vd1_axi_arprot,
    output wire [3:0]               s02_vd1_axi_arqos,
    output wire [3:0]               s02_vd1_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s02_vd1_axi_aruser,
    output wire                     s02_vd1_axi_arvalid,
    input  wire                     s02_vd1_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd1_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s02_vd1_axi_rdata,
    input  wire [1:0]               s02_vd1_axi_rresp,
    input  wire                     s02_vd1_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s02_vd1_axi_ruser,
    input  wire                     s02_vd1_axi_rvalid,
    output wire                     s02_vd1_axi_rready,
//vd2
    output wire [M_ID_WIDTH-1:0]    s00_vd2_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s00_vd2_axi_awaddr,
    output wire [7:0]               s00_vd2_axi_awlen,
    output wire [2:0]               s00_vd2_axi_awsize,
    output wire [1:0]               s00_vd2_axi_awburst,
    output wire                     s00_vd2_axi_awlock,
    output wire [3:0]               s00_vd2_axi_awcache,
    output wire [2:0]               s00_vd2_axi_awprot,
    output wire [3:0]               s00_vd2_axi_awqos,
    output wire [3:0]               s00_vd2_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s00_vd2_axi_awuser,
    output wire                     s00_vd2_axi_awvalid,
    input  wire                     s00_vd2_axi_awready,
    output wire [DATA_WIDTH-1:0]    s00_vd2_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s00_vd2_axi_wstrb,
    output wire                     s00_vd2_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s00_vd2_axi_wuser,
    output wire                     s00_vd2_axi_wvalid,
    input  wire                     s00_vd2_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd2_axi_bid,
    input  wire [1:0]               s00_vd2_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s00_vd2_axi_buser,
    input  wire                     s00_vd2_axi_bvalid,
    output wire                     s00_vd2_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s00_vd2_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s00_vd2_axi_araddr,
    output wire [7:0]               s00_vd2_axi_arlen,
    output wire [2:0]               s00_vd2_axi_arsize,
    output wire [1:0]               s00_vd2_axi_arburst,
    output wire                     s00_vd2_axi_arlock,
    output wire [3:0]               s00_vd2_axi_arcache,
    output wire [2:0]               s00_vd2_axi_arprot,
    output wire [3:0]               s00_vd2_axi_arqos,
    output wire [3:0]               s00_vd2_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s00_vd2_axi_aruser,
    output wire                     s00_vd2_axi_arvalid,
    input  wire                     s00_vd2_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd2_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s00_vd2_axi_rdata,
    input  wire [1:0]               s00_vd2_axi_rresp,
    input  wire                     s00_vd2_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s00_vd2_axi_ruser,
    input  wire                     s00_vd2_axi_rvalid,
    output wire                     s00_vd2_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s01_vd2_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s01_vd2_axi_awaddr,
    output wire [7:0]               s01_vd2_axi_awlen,
    output wire [2:0]               s01_vd2_axi_awsize,
    output wire [1:0]               s01_vd2_axi_awburst,
    output wire                     s01_vd2_axi_awlock,
    output wire [3:0]               s01_vd2_axi_awcache,
    output wire [2:0]               s01_vd2_axi_awprot,
    output wire [3:0]               s01_vd2_axi_awqos,
    output wire [3:0]               s01_vd2_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s01_vd2_axi_awuser,
    output wire                     s01_vd2_axi_awvalid,
    input  wire                     s01_vd2_axi_awready,
    output wire [DATA_WIDTH-1:0]    s01_vd2_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s01_vd2_axi_wstrb,
    output wire                     s01_vd2_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s01_vd2_axi_wuser,
    output wire                     s01_vd2_axi_wvalid,
    input  wire                     s01_vd2_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd2_axi_bid,
    input  wire [1:0]               s01_vd2_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s01_vd2_axi_buser,
    input  wire                     s01_vd2_axi_bvalid,
    output wire                     s01_vd2_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s01_vd2_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s01_vd2_axi_araddr,
    output wire [7:0]               s01_vd2_axi_arlen,
    output wire [2:0]               s01_vd2_axi_arsize,
    output wire [1:0]               s01_vd2_axi_arburst,
    output wire                     s01_vd2_axi_arlock,
    output wire [3:0]               s01_vd2_axi_arcache,
    output wire [2:0]               s01_vd2_axi_arprot,
    output wire [3:0]               s01_vd2_axi_arqos,
    output wire [3:0]               s01_vd2_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s01_vd2_axi_aruser,
    output wire                     s01_vd2_axi_arvalid,
    input  wire                     s01_vd2_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd2_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s01_vd2_axi_rdata,
    input  wire [1:0]               s01_vd2_axi_rresp,
    input  wire                     s01_vd2_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s01_vd2_axi_ruser,
    input  wire                     s01_vd2_axi_rvalid,
    output wire                     s01_vd2_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s02_vd2_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s02_vd2_axi_awaddr,
    output wire [7:0]               s02_vd2_axi_awlen,
    output wire [2:0]               s02_vd2_axi_awsize,
    output wire [1:0]               s02_vd2_axi_awburst,
    output wire                     s02_vd2_axi_awlock,
    output wire [3:0]               s02_vd2_axi_awcache,
    output wire [2:0]               s02_vd2_axi_awprot,
    output wire [3:0]               s02_vd2_axi_awqos,
    output wire [3:0]               s02_vd2_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s02_vd2_axi_awuser,
    output wire                     s02_vd2_axi_awvalid,
    input  wire                     s02_vd2_axi_awready,
    output wire [DATA_WIDTH-1:0]    s02_vd2_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s02_vd2_axi_wstrb,
    output wire                     s02_vd2_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s02_vd2_axi_wuser,
    output wire                     s02_vd2_axi_wvalid,
    input  wire                     s02_vd2_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd2_axi_bid,
    input  wire [1:0]               s02_vd2_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s02_vd2_axi_buser,
    input  wire                     s02_vd2_axi_bvalid,
    output wire                     s02_vd2_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s02_vd2_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s02_vd2_axi_araddr,
    output wire [7:0]               s02_vd2_axi_arlen,
    output wire [2:0]               s02_vd2_axi_arsize,
    output wire [1:0]               s02_vd2_axi_arburst,
    output wire                     s02_vd2_axi_arlock,
    output wire [3:0]               s02_vd2_axi_arcache,
    output wire [2:0]               s02_vd2_axi_arprot,
    output wire [3:0]               s02_vd2_axi_arqos,
    output wire [3:0]               s02_vd2_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s02_vd2_axi_aruser,
    output wire                     s02_vd2_axi_arvalid,
    input  wire                     s02_vd2_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd2_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s02_vd2_axi_rdata,
    input  wire [1:0]               s02_vd2_axi_rresp,
    input  wire                     s02_vd2_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s02_vd2_axi_ruser,
    input  wire                     s02_vd2_axi_rvalid,
    output wire                     s02_vd2_axi_rready,
//vd3
    output wire [M_ID_WIDTH-1:0]    s00_vd3_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s00_vd3_axi_awaddr,
    output wire [7:0]               s00_vd3_axi_awlen,
    output wire [2:0]               s00_vd3_axi_awsize,
    output wire [1:0]               s00_vd3_axi_awburst,
    output wire                     s00_vd3_axi_awlock,
    output wire [3:0]               s00_vd3_axi_awcache,
    output wire [2:0]               s00_vd3_axi_awprot,
    output wire [3:0]               s00_vd3_axi_awqos,
    output wire [3:0]               s00_vd3_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s00_vd3_axi_awuser,
    output wire                     s00_vd3_axi_awvalid,
    input  wire                     s00_vd3_axi_awready,
    output wire [DATA_WIDTH-1:0]    s00_vd3_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s00_vd3_axi_wstrb,
    output wire                     s00_vd3_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s00_vd3_axi_wuser,
    output wire                     s00_vd3_axi_wvalid,
    input  wire                     s00_vd3_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd3_axi_bid,
    input  wire [1:0]               s00_vd3_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s00_vd3_axi_buser,
    input  wire                     s00_vd3_axi_bvalid,
    output wire                     s00_vd3_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s00_vd3_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s00_vd3_axi_araddr,
    output wire [7:0]               s00_vd3_axi_arlen,
    output wire [2:0]               s00_vd3_axi_arsize,
    output wire [1:0]               s00_vd3_axi_arburst,
    output wire                     s00_vd3_axi_arlock,
    output wire [3:0]               s00_vd3_axi_arcache,
    output wire [2:0]               s00_vd3_axi_arprot,
    output wire [3:0]               s00_vd3_axi_arqos,
    output wire [3:0]               s00_vd3_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s00_vd3_axi_aruser,
    output wire                     s00_vd3_axi_arvalid,
    input  wire                     s00_vd3_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s00_vd3_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s00_vd3_axi_rdata,
    input  wire [1:0]               s00_vd3_axi_rresp,
    input  wire                     s00_vd3_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s00_vd3_axi_ruser,
    input  wire                     s00_vd3_axi_rvalid,
    output wire                     s00_vd3_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s01_vd3_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s01_vd3_axi_awaddr,
    output wire [7:0]               s01_vd3_axi_awlen,
    output wire [2:0]               s01_vd3_axi_awsize,
    output wire [1:0]               s01_vd3_axi_awburst,
    output wire                     s01_vd3_axi_awlock,
    output wire [3:0]               s01_vd3_axi_awcache,
    output wire [2:0]               s01_vd3_axi_awprot,
    output wire [3:0]               s01_vd3_axi_awqos,
    output wire [3:0]               s01_vd3_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s01_vd3_axi_awuser,
    output wire                     s01_vd3_axi_awvalid,
    input  wire                     s01_vd3_axi_awready,
    output wire [DATA_WIDTH-1:0]    s01_vd3_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s01_vd3_axi_wstrb,
    output wire                     s01_vd3_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s01_vd3_axi_wuser,
    output wire                     s01_vd3_axi_wvalid,
    input  wire                     s01_vd3_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd3_axi_bid,
    input  wire [1:0]               s01_vd3_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s01_vd3_axi_buser,
    input  wire                     s01_vd3_axi_bvalid,
    output wire                     s01_vd3_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s01_vd3_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s01_vd3_axi_araddr,
    output wire [7:0]               s01_vd3_axi_arlen,
    output wire [2:0]               s01_vd3_axi_arsize,
    output wire [1:0]               s01_vd3_axi_arburst,
    output wire                     s01_vd3_axi_arlock,
    output wire [3:0]               s01_vd3_axi_arcache,
    output wire [2:0]               s01_vd3_axi_arprot,
    output wire [3:0]               s01_vd3_axi_arqos,
    output wire [3:0]               s01_vd3_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s01_vd3_axi_aruser,
    output wire                     s01_vd3_axi_arvalid,
    input  wire                     s01_vd3_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s01_vd3_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s01_vd3_axi_rdata,
    input  wire [1:0]               s01_vd3_axi_rresp,
    input  wire                     s01_vd3_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s01_vd3_axi_ruser,
    input  wire                     s01_vd3_axi_rvalid,
    output wire                     s01_vd3_axi_rready,

    output wire [M_ID_WIDTH-1:0]    s02_vd3_axi_awid,
    output wire [ADDR_WIDTH-1:0]    s02_vd3_axi_awaddr,
    output wire [7:0]               s02_vd3_axi_awlen,
    output wire [2:0]               s02_vd3_axi_awsize,
    output wire [1:0]               s02_vd3_axi_awburst,
    output wire                     s02_vd3_axi_awlock,
    output wire [3:0]               s02_vd3_axi_awcache,
    output wire [2:0]               s02_vd3_axi_awprot,
    output wire [3:0]               s02_vd3_axi_awqos,
    output wire [3:0]               s02_vd3_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  s02_vd3_axi_awuser,
    output wire                     s02_vd3_axi_awvalid,
    input  wire                     s02_vd3_axi_awready,
    output wire [DATA_WIDTH-1:0]    s02_vd3_axi_wdata,
    output wire [STRB_WIDTH-1:0]    s02_vd3_axi_wstrb,
    output wire                     s02_vd3_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   s02_vd3_axi_wuser,
    output wire                     s02_vd3_axi_wvalid,
    input  wire                     s02_vd3_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd3_axi_bid,
    input  wire [1:0]               s02_vd3_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   s02_vd3_axi_buser,
    input  wire                     s02_vd3_axi_bvalid,
    output wire                     s02_vd3_axi_bready,
    output wire [M_ID_WIDTH-1:0]    s02_vd3_axi_arid,
    output wire [ADDR_WIDTH-1:0]    s02_vd3_axi_araddr,
    output wire [7:0]               s02_vd3_axi_arlen,
    output wire [2:0]               s02_vd3_axi_arsize,
    output wire [1:0]               s02_vd3_axi_arburst,
    output wire                     s02_vd3_axi_arlock,
    output wire [3:0]               s02_vd3_axi_arcache,
    output wire [2:0]               s02_vd3_axi_arprot,
    output wire [3:0]               s02_vd3_axi_arqos,
    output wire [3:0]               s02_vd3_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  s02_vd3_axi_aruser,
    output wire                     s02_vd3_axi_arvalid,
    input  wire                     s02_vd3_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    s02_vd3_axi_rid,
    input  wire [DATA_WIDTH-1:0]    s02_vd3_axi_rdata,
    input  wire [1:0]               s02_vd3_axi_rresp,
    input  wire                     s02_vd3_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   s02_vd3_axi_ruser,
    input  wire                     s02_vd3_axi_rvalid,
    output wire                     s02_vd3_axi_rready,
/* AXI master interface
*/
    output wire [M_ID_WIDTH-1:0]    m00_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m00_axi_awaddr,
    output wire [7:0]               m00_axi_awlen,
    output wire [2:0]               m00_axi_awsize,
    output wire [1:0]               m00_axi_awburst,
    output wire                     m00_axi_awlock,
    output wire [3:0]               m00_axi_awcache,
    output wire [2:0]               m00_axi_awprot,
    output wire [3:0]               m00_axi_awqos,
    output wire [3:0]               m00_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m00_axi_awuser,
    output wire                     m00_axi_awvalid,
    input  wire                     m00_axi_awready,
    output wire [DATA_WIDTH-1:0]    m00_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m00_axi_wstrb,
    output wire                     m00_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m00_axi_wuser,
    output wire                     m00_axi_wvalid,
    input  wire                     m00_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    m00_axi_bid,
    input  wire [1:0]               m00_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m00_axi_buser,
    input  wire                     m00_axi_bvalid,
    output wire                     m00_axi_bready,
    output wire [M_ID_WIDTH-1:0]    m00_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m00_axi_araddr,
    output wire [7:0]               m00_axi_arlen,
    output wire [2:0]               m00_axi_arsize,
    output wire [1:0]               m00_axi_arburst,
    output wire                     m00_axi_arlock,
    output wire [3:0]               m00_axi_arcache,
    output wire [2:0]               m00_axi_arprot,
    output wire [3:0]               m00_axi_arqos,
    output wire [3:0]               m00_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m00_axi_aruser,
    output wire                     m00_axi_arvalid,
    input  wire                     m00_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    m00_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m00_axi_rdata,
    input  wire [1:0]               m00_axi_rresp,
    input  wire                     m00_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m00_axi_ruser,
    input  wire                     m00_axi_rvalid,
    output wire                     m00_axi_rready,

    output wire [M_ID_WIDTH-1:0]    m01_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m01_axi_awaddr,
    output wire [7:0]               m01_axi_awlen,
    output wire [2:0]               m01_axi_awsize,
    output wire [1:0]               m01_axi_awburst,
    output wire                     m01_axi_awlock,
    output wire [3:0]               m01_axi_awcache,
    output wire [2:0]               m01_axi_awprot,
    output wire [3:0]               m01_axi_awqos,
    output wire [3:0]               m01_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m01_axi_awuser,
    output wire                     m01_axi_awvalid,
    input  wire                     m01_axi_awready,
    output wire [DATA_WIDTH-1:0]    m01_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m01_axi_wstrb,
    output wire                     m01_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m01_axi_wuser,
    output wire                     m01_axi_wvalid,
    input  wire                     m01_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    m01_axi_bid,
    input  wire [1:0]               m01_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m01_axi_buser,
    input  wire                     m01_axi_bvalid,
    output wire                     m01_axi_bready,
    output wire [M_ID_WIDTH-1:0]    m01_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m01_axi_araddr,
    output wire [7:0]               m01_axi_arlen,
    output wire [2:0]               m01_axi_arsize,
    output wire [1:0]               m01_axi_arburst,
    output wire                     m01_axi_arlock,
    output wire [3:0]               m01_axi_arcache,
    output wire [2:0]               m01_axi_arprot,
    output wire [3:0]               m01_axi_arqos,
    output wire [3:0]               m01_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m01_axi_aruser,
    output wire                     m01_axi_arvalid,
    input  wire                     m01_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    m01_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m01_axi_rdata,
    input  wire [1:0]               m01_axi_rresp,
    input  wire                     m01_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m01_axi_ruser,
    input  wire                     m01_axi_rvalid,
    output wire                     m01_axi_rready,

    output wire [M_ID_WIDTH-1:0]    m02_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m02_axi_awaddr,
    output wire [7:0]               m02_axi_awlen,
    output wire [2:0]               m02_axi_awsize,
    output wire [1:0]               m02_axi_awburst,
    output wire                     m02_axi_awlock,
    output wire [3:0]               m02_axi_awcache,
    output wire [2:0]               m02_axi_awprot,
    output wire [3:0]               m02_axi_awqos,
    output wire [3:0]               m02_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m02_axi_awuser,
    output wire                     m02_axi_awvalid,
    input  wire                     m02_axi_awready,
    output wire [DATA_WIDTH-1:0]    m02_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m02_axi_wstrb,
    output wire                     m02_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m02_axi_wuser,
    output wire                     m02_axi_wvalid,
    input  wire                     m02_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    m02_axi_bid,
    input  wire [1:0]               m02_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m02_axi_buser,
    input  wire                     m02_axi_bvalid,
    output wire                     m02_axi_bready,
    output wire [M_ID_WIDTH-1:0]    m02_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m02_axi_araddr,
    output wire [7:0]               m02_axi_arlen,
    output wire [2:0]               m02_axi_arsize,
    output wire [1:0]               m02_axi_arburst,
    output wire                     m02_axi_arlock,
    output wire [3:0]               m02_axi_arcache,
    output wire [2:0]               m02_axi_arprot,
    output wire [3:0]               m02_axi_arqos,
    output wire [3:0]               m02_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m02_axi_aruser,
    output wire                     m02_axi_arvalid,
    input  wire                     m02_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    m02_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m02_axi_rdata,
    input  wire [1:0]               m02_axi_rresp,
    input  wire                     m02_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m02_axi_ruser,
    input  wire                     m02_axi_rvalid,
    output wire                     m02_axi_rready,

    output wire [M_ID_WIDTH-1:0]    m03_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m03_axi_awaddr,
    output wire [7:0]               m03_axi_awlen,
    output wire [2:0]               m03_axi_awsize,
    output wire [1:0]               m03_axi_awburst,
    output wire                     m03_axi_awlock,
    output wire [3:0]               m03_axi_awcache,
    output wire [2:0]               m03_axi_awprot,
    output wire [3:0]               m03_axi_awqos,
    output wire [3:0]               m03_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m03_axi_awuser,
    output wire                     m03_axi_awvalid,
    input  wire                     m03_axi_awready,
    output wire [DATA_WIDTH-1:0]    m03_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m03_axi_wstrb,
    output wire                     m03_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m03_axi_wuser,
    output wire                     m03_axi_wvalid,
    input  wire                     m03_axi_wready,
    input  wire [M_ID_WIDTH-1:0]    m03_axi_bid,
    input  wire [1:0]               m03_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m03_axi_buser,
    input  wire                     m03_axi_bvalid,
    output wire                     m03_axi_bready,
    output wire [M_ID_WIDTH-1:0]    m03_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m03_axi_araddr,
    output wire [7:0]               m03_axi_arlen,
    output wire [2:0]               m03_axi_arsize,
    output wire [1:0]               m03_axi_arburst,
    output wire                     m03_axi_arlock,
    output wire [3:0]               m03_axi_arcache,
    output wire [2:0]               m03_axi_arprot,
    output wire [3:0]               m03_axi_arqos,
    output wire [3:0]               m03_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m03_axi_aruser,
    output wire                     m03_axi_arvalid,
    input  wire                     m03_axi_arready,
    input  wire [M_ID_WIDTH-1:0]    m03_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m03_axi_rdata,
    input  wire [1:0]               m03_axi_rresp,
    input  wire                     m03_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m03_axi_ruser,
    input  wire                     m03_axi_rvalid,
    output wire                     m03_axi_rready
);

//inst0
//m00+vd0
axi_tmr_voter_ds_1m3s#(
   .DATA_WIDTH     (64             ),
   .ADDR_WIDTH     (32             ),
   .STRB_WIDTH     ((DATA_WIDTH/8) ),
   .S_ID_WIDTH     (8              ),
   .M_ID_WIDTH     (S_ID_WIDTH+$clog2(3)),
   .AWUSER_ENABLE  (0              ),
   .AWUSER_WIDTH   (1              ),
   .WUSER_ENABLE   (0              ),
   .WUSER_WIDTH    (1              ),
   .BUSER_ENABLE   (0              ),
   .BUSER_WIDTH    (1              ),
   .ARUSER_ENABLE  (0              ),
   .ARUSER_WIDTH   (1              ),
   .RUSER_ENABLE   (0              ),
   .RUSER_WIDTH    (1              ),
   .S00_THREADS    (8              ),
   .S00_ACCEPT     (16             ),
   .S01_THREADS    (8              ),
   .S01_ACCEPT     (16             ),
   .S02_THREADS    (8              ),
   .S02_ACCEPT     (16             ),
   .M_REGIONS      (1              ),
   .M00_BASE_ADDR  (0              ),
   .M00_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M00_CONNECT_READ(3'b100         ),
   .M00_CONNECT_WRITE(3'b100         ),
   .M00_ISSUE      (8              ),
   .M00_SECURE     (1              ),
   .M01_BASE_ADDR  (0              ),
   .M01_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M01_CONNECT_READ(3'b011         ),
   .M01_CONNECT_WRITE(3'b011         ),
   .M01_ISSUE      (8              ),
   .M01_SECURE     (0              ),
   .M02_BASE_ADDR  (0              ),
   .M02_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M02_CONNECT_READ(3'b100         ),
   .M02_CONNECT_WRITE(3'b100         ),
   .M02_ISSUE      (8              ),
   .M02_SECURE     (1              ),
   .M03_BASE_ADDR  (0              ),
   .M03_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M03_CONNECT_READ(3'b011         ),
   .M03_CONNECT_WRITE(3'b011         ),
   .M03_ISSUE      (8              ),
   .M03_SECURE     (0              ),
   .S00_AW_REG_TYPE(0              ),
   .S00_W_REG_TYPE (0              ),
   .S00_B_REG_TYPE (1              ),
   .S00_AR_REG_TYPE(0              ),
   .S00_R_REG_TYPE (2              ),
   .S01_AW_REG_TYPE(0              ),
   .S01_W_REG_TYPE (0              ),
   .S01_B_REG_TYPE (1              ),
   .S01_AR_REG_TYPE(0              ),
   .S01_R_REG_TYPE (2              ),
   .S02_AW_REG_TYPE(0              ),
   .S02_W_REG_TYPE (0              ),
   .S02_B_REG_TYPE (1              ),
   .S02_AR_REG_TYPE(0              ),
   .S02_R_REG_TYPE (2              ),
   .M00_AW_REG_TYPE(1              ),
   .M00_W_REG_TYPE (2              ),
   .M00_B_REG_TYPE (0              ),
   .M00_AR_REG_TYPE(1              ),
   .M00_R_REG_TYPE (0              ),
   .M01_AW_REG_TYPE(1              ),
   .M01_W_REG_TYPE (2              ),
   .M01_B_REG_TYPE (0              ),
   .M01_AR_REG_TYPE(1              ),
   .M01_R_REG_TYPE (0              ),
   .M02_AW_REG_TYPE(1              ),
   .M02_W_REG_TYPE (2              ),
   .M02_B_REG_TYPE (0              ),
   .M02_AR_REG_TYPE(1              ),
   .M02_R_REG_TYPE (0              ),
   .M03_AW_REG_TYPE(1              ),
   .M03_W_REG_TYPE (2              ),
   .M03_B_REG_TYPE (0              ),
   .M03_AR_REG_TYPE(1              ),
   .M03_R_REG_TYPE (0              )
)
 u_axi_tmr_voter_ds_1m3s_inst0(
    .clk                                (clk                       ),
    .rst                                (rst                       ),
//s00
    .s00_axi_awid                       (s00_vd0_axi_awid              ),
    .s00_axi_awaddr                     (s00_vd0_axi_awaddr            ),
    .s00_axi_awlen                      (s00_vd0_axi_awlen             ),
    .s00_axi_awsize                     (s00_vd0_axi_awsize            ),
    .s00_axi_awburst                    (s00_vd0_axi_awburst           ),
    .s00_axi_awlock                     (s00_vd0_axi_awlock            ),
    .s00_axi_awcache                    (s00_vd0_axi_awcache           ),
    .s00_axi_awprot                     (s00_vd0_axi_awprot            ),
    .s00_axi_awqos                      (s00_vd0_axi_awqos             ),
    .s00_axi_awregion                   (s00_vd0_axi_awregion          ),
    .s00_axi_awuser                     (s00_vd0_axi_awuser            ),
    .s00_axi_awvalid                    (s00_vd0_axi_awvalid           ),
    .s00_axi_awready                    (s00_vd0_axi_awready           ),
    .s00_axi_wdata                      (s00_vd0_axi_wdata             ),
    .s00_axi_wstrb                      (s00_vd0_axi_wstrb             ),
    .s00_axi_wlast                      (s00_vd0_axi_wlast             ),
    .s00_axi_wuser                      (s00_vd0_axi_wuser             ),
    .s00_axi_wvalid                     (s00_vd0_axi_wvalid            ),
    .s00_axi_wready                     (s00_vd0_axi_wready            ),
    .s00_axi_bid                        (s00_vd0_axi_bid               ),
    .s00_axi_bresp                      (s00_vd0_axi_bresp             ),
    .s00_axi_buser                      (s00_vd0_axi_buser             ),
    .s00_axi_bvalid                     (s00_vd0_axi_bvalid            ),
    .s00_axi_bready                     (s00_vd0_axi_bready            ),
    .s00_axi_arid                       (s00_vd0_axi_arid              ),
    .s00_axi_araddr                     (s00_vd0_axi_araddr            ),
    .s00_axi_arlen                      (s00_vd0_axi_arlen             ),
    .s00_axi_arsize                     (s00_vd0_axi_arsize            ),
    .s00_axi_arburst                    (s00_vd0_axi_arburst           ),
    .s00_axi_arlock                     (s00_vd0_axi_arlock            ),
    .s00_axi_arcache                    (s00_vd0_axi_arcache           ),
    .s00_axi_arprot                     (s00_vd0_axi_arprot            ),
    .s00_axi_arqos                      (s00_vd0_axi_arqos             ),
    .s00_axi_arregion                   (s00_vd0_axi_arregion          ),
    .s00_axi_aruser                     (s00_vd0_axi_aruser            ),
    .s00_axi_arvalid                    (s00_vd0_axi_arvalid           ),
    .s00_axi_arready                    (s00_vd0_axi_arready           ),
    .s00_axi_rid                        (s00_vd0_axi_rid               ),
    .s00_axi_rdata                      (s00_vd0_axi_rdata             ),
    .s00_axi_rresp                      (s00_vd0_axi_rresp             ),
    .s00_axi_rlast                      (s00_vd0_axi_rlast             ),
    .s00_axi_ruser                      (s00_vd0_axi_ruser             ),
    .s00_axi_rvalid                     (s00_vd0_axi_rvalid            ),
    .s00_axi_rready                     (s00_vd0_axi_rready            ),
//s01
    .s01_axi_awid                       (s01_vd0_axi_awid              ),
    .s01_axi_awaddr                     (s01_vd0_axi_awaddr            ),
    .s01_axi_awlen                      (s01_vd0_axi_awlen             ),
    .s01_axi_awsize                     (s01_vd0_axi_awsize            ),
    .s01_axi_awburst                    (s01_vd0_axi_awburst           ),
    .s01_axi_awlock                     (s01_vd0_axi_awlock            ),
    .s01_axi_awcache                    (s01_vd0_axi_awcache           ),
    .s01_axi_awprot                     (s01_vd0_axi_awprot            ),
    .s01_axi_awqos                      (s01_vd0_axi_awqos             ),
    .s01_axi_awregion                   (s01_vd0_axi_awregion          ),
    .s01_axi_awuser                     (s01_vd0_axi_awuser            ),
    .s01_axi_awvalid                    (s01_vd0_axi_awvalid           ),
    .s01_axi_awready                    (s01_vd0_axi_awready           ),
    .s01_axi_wdata                      (s01_vd0_axi_wdata             ),
    .s01_axi_wstrb                      (s01_vd0_axi_wstrb             ),
    .s01_axi_wlast                      (s01_vd0_axi_wlast             ),
    .s01_axi_wuser                      (s01_vd0_axi_wuser             ),
    .s01_axi_wvalid                     (s01_vd0_axi_wvalid            ),
    .s01_axi_wready                     (s01_vd0_axi_wready            ),
    .s01_axi_bid                        (s01_vd0_axi_bid               ),
    .s01_axi_bresp                      (s01_vd0_axi_bresp             ),
    .s01_axi_buser                      (s01_vd0_axi_buser             ),
    .s01_axi_bvalid                     (s01_vd0_axi_bvalid            ),
    .s01_axi_bready                     (s01_vd0_axi_bready            ),
    .s01_axi_arid                       (s01_vd0_axi_arid              ),
    .s01_axi_araddr                     (s01_vd0_axi_araddr            ),
    .s01_axi_arlen                      (s01_vd0_axi_arlen             ),
    .s01_axi_arsize                     (s01_vd0_axi_arsize            ),
    .s01_axi_arburst                    (s01_vd0_axi_arburst           ),
    .s01_axi_arlock                     (s01_vd0_axi_arlock            ),
    .s01_axi_arcache                    (s01_vd0_axi_arcache           ),
    .s01_axi_arprot                     (s01_vd0_axi_arprot            ),
    .s01_axi_arqos                      (s01_vd0_axi_arqos             ),
    .s01_axi_arregion                   (s01_vd0_axi_arregion          ),
    .s01_axi_aruser                     (s01_vd0_axi_aruser            ),
    .s01_axi_arvalid                    (s01_vd0_axi_arvalid           ),
    .s01_axi_arready                    (s01_vd0_axi_arready           ),
    .s01_axi_rid                        (s01_vd0_axi_rid               ),
    .s01_axi_rdata                      (s01_vd0_axi_rdata             ),
    .s01_axi_rresp                      (s01_vd0_axi_rresp             ),
    .s01_axi_rlast                      (s01_vd0_axi_rlast             ),
    .s01_axi_ruser                      (s01_vd0_axi_ruser             ),
    .s01_axi_rvalid                     (s01_vd0_axi_rvalid            ),
    .s01_axi_rready                     (s01_vd0_axi_rready            ),
//s02
    .s02_axi_awid                       (s02_vd0_axi_awid              ),
    .s02_axi_awaddr                     (s02_vd0_axi_awaddr            ),
    .s02_axi_awlen                      (s02_vd0_axi_awlen             ),
    .s02_axi_awsize                     (s02_vd0_axi_awsize            ),
    .s02_axi_awburst                    (s02_vd0_axi_awburst           ),
    .s02_axi_awlock                     (s02_vd0_axi_awlock            ),
    .s02_axi_awcache                    (s02_vd0_axi_awcache           ),
    .s02_axi_awprot                     (s02_vd0_axi_awprot            ),
    .s02_axi_awqos                      (s02_vd0_axi_awqos             ),
    .s02_axi_awregion                   (s02_vd0_axi_awregion          ),
    .s02_axi_awuser                     (s02_vd0_axi_awuser            ),
    .s02_axi_awvalid                    (s02_vd0_axi_awvalid           ),
    .s02_axi_awready                    (s02_vd0_axi_awready           ),
    .s02_axi_wdata                      (s02_vd0_axi_wdata             ),
    .s02_axi_wstrb                      (s02_vd0_axi_wstrb             ),
    .s02_axi_wlast                      (s02_vd0_axi_wlast             ),
    .s02_axi_wuser                      (s02_vd0_axi_wuser             ),
    .s02_axi_wvalid                     (s02_vd0_axi_wvalid            ),
    .s02_axi_wready                     (s02_vd0_axi_wready            ),
    .s02_axi_bid                        (s02_vd0_axi_bid               ),
    .s02_axi_bresp                      (s02_vd0_axi_bresp             ),
    .s02_axi_buser                      (s02_vd0_axi_buser             ),
    .s02_axi_bvalid                     (s02_vd0_axi_bvalid            ),
    .s02_axi_bready                     (s02_vd0_axi_bready            ),
    .s02_axi_arid                       (s02_vd0_axi_arid              ),
    .s02_axi_araddr                     (s02_vd0_axi_araddr            ),
    .s02_axi_arlen                      (s02_vd0_axi_arlen             ),
    .s02_axi_arsize                     (s02_vd0_axi_arsize            ),
    .s02_axi_arburst                    (s02_vd0_axi_arburst           ),
    .s02_axi_arlock                     (s02_vd0_axi_arlock            ),
    .s02_axi_arcache                    (s02_vd0_axi_arcache           ),
    .s02_axi_arprot                     (s02_vd0_axi_arprot            ),
    .s02_axi_arqos                      (s02_vd0_axi_arqos             ),
    .s02_axi_arregion                   (s02_vd0_axi_arregion          ),
    .s02_axi_aruser                     (s02_vd0_axi_aruser            ),
    .s02_axi_arvalid                    (s02_vd0_axi_arvalid           ),
    .s02_axi_arready                    (s02_vd0_axi_arready           ),
    .s02_axi_rid                        (s02_vd0_axi_rid               ),
    .s02_axi_rdata                      (s02_vd0_axi_rdata             ),
    .s02_axi_rresp                      (s02_vd0_axi_rresp             ),
    .s02_axi_rlast                      (s02_vd0_axi_rlast             ),
    .s02_axi_ruser                      (s02_vd0_axi_ruser             ),
    .s02_axi_rvalid                     (s02_vd0_axi_rvalid            ),
    .s02_axi_rready                     (s02_vd0_axi_rready            ),
//m00
    .m00_axi_awid                       (m00_axi_awid              ),
    .m00_axi_awaddr                     (m00_axi_awaddr            ),
    .m00_axi_awlen                      (m00_axi_awlen             ),
    .m00_axi_awsize                     (m00_axi_awsize            ),
    .m00_axi_awburst                    (m00_axi_awburst           ),
    .m00_axi_awlock                     (m00_axi_awlock            ),
    .m00_axi_awcache                    (m00_axi_awcache           ),
    .m00_axi_awprot                     (m00_axi_awprot            ),
    .m00_axi_awqos                      (m00_axi_awqos             ),
    .m00_axi_awregion                   (m00_axi_awregion          ),
    .m00_axi_awuser                     (m00_axi_awuser            ),
    .m00_axi_awvalid                    (m00_axi_awvalid           ),
    .m00_axi_awready                    (m00_axi_awready           ),
    .m00_axi_wdata                      (m00_axi_wdata             ),
    .m00_axi_wstrb                      (m00_axi_wstrb             ),
    .m00_axi_wlast                      (m00_axi_wlast             ),
    .m00_axi_wuser                      (m00_axi_wuser             ),
    .m00_axi_wvalid                     (m00_axi_wvalid            ),
    .m00_axi_wready                     (m00_axi_wready            ),
    .m00_axi_bid                        (m00_axi_bid               ),
    .m00_axi_bresp                      (m00_axi_bresp             ),
    .m00_axi_buser                      (m00_axi_buser             ),
    .m00_axi_bvalid                     (m00_axi_bvalid            ),
    .m00_axi_bready                     (m00_axi_bready            ),
    .m00_axi_arid                       (m00_axi_arid              ),
    .m00_axi_araddr                     (m00_axi_araddr            ),
    .m00_axi_arlen                      (m00_axi_arlen             ),
    .m00_axi_arsize                     (m00_axi_arsize            ),
    .m00_axi_arburst                    (m00_axi_arburst           ),
    .m00_axi_arlock                     (m00_axi_arlock            ),
    .m00_axi_arcache                    (m00_axi_arcache           ),
    .m00_axi_arprot                     (m00_axi_arprot            ),
    .m00_axi_arqos                      (m00_axi_arqos             ),
    .m00_axi_arregion                   (m00_axi_arregion          ),
    .m00_axi_aruser                     (m00_axi_aruser            ),
    .m00_axi_arvalid                    (m00_axi_arvalid           ),
    .m00_axi_arready                    (m00_axi_arready           ),
    .m00_axi_rid                        (m00_axi_rid               ),
    .m00_axi_rdata                      (m00_axi_rdata             ),
    .m00_axi_rresp                      (m00_axi_rresp             ),
    .m00_axi_rlast                      (m00_axi_rlast             ),
    .m00_axi_ruser                      (m00_axi_ruser             ),
    .m00_axi_rvalid                     (m00_axi_rvalid            ),
    .m00_axi_rready                     (m00_axi_rready            )
);

//inst1
//m01+vd1
axi_tmr_voter_ds_1m3s#(
   .DATA_WIDTH     (64             ),
   .ADDR_WIDTH     (32             ),
   .STRB_WIDTH     ((DATA_WIDTH/8) ),
   .S_ID_WIDTH     (8              ),
   .M_ID_WIDTH     (S_ID_WIDTH+$clog2(3)),
   .AWUSER_ENABLE  (0              ),
   .AWUSER_WIDTH   (1              ),
   .WUSER_ENABLE   (0              ),
   .WUSER_WIDTH    (1              ),
   .BUSER_ENABLE   (0              ),
   .BUSER_WIDTH    (1              ),
   .ARUSER_ENABLE  (0              ),
   .ARUSER_WIDTH   (1              ),
   .RUSER_ENABLE   (0              ),
   .RUSER_WIDTH    (1              ),
   .S00_THREADS    (8              ),
   .S00_ACCEPT     (16             ),
   .S01_THREADS    (8              ),
   .S01_ACCEPT     (16             ),
   .S02_THREADS    (8              ),
   .S02_ACCEPT     (16             ),
   .M_REGIONS      (1              ),
   .M00_BASE_ADDR  (0              ),
   .M00_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M00_CONNECT_READ(3'b100         ),
   .M00_CONNECT_WRITE(3'b100         ),
   .M00_ISSUE      (8              ),
   .M00_SECURE     (1              ),
   .M01_BASE_ADDR  (0              ),
   .M01_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M01_CONNECT_READ(3'b011         ),
   .M01_CONNECT_WRITE(3'b011         ),
   .M01_ISSUE      (8              ),
   .M01_SECURE     (0              ),
   .M02_BASE_ADDR  (0              ),
   .M02_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M02_CONNECT_READ(3'b100         ),
   .M02_CONNECT_WRITE(3'b100         ),
   .M02_ISSUE      (8              ),
   .M02_SECURE     (1              ),
   .M03_BASE_ADDR  (0              ),
   .M03_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M03_CONNECT_READ(3'b011         ),
   .M03_CONNECT_WRITE(3'b011         ),
   .M03_ISSUE      (8              ),
   .M03_SECURE     (0              ),
   .S00_AW_REG_TYPE(0              ),
   .S00_W_REG_TYPE (0              ),
   .S00_B_REG_TYPE (1              ),
   .S00_AR_REG_TYPE(0              ),
   .S00_R_REG_TYPE (2              ),
   .S01_AW_REG_TYPE(0              ),
   .S01_W_REG_TYPE (0              ),
   .S01_B_REG_TYPE (1              ),
   .S01_AR_REG_TYPE(0              ),
   .S01_R_REG_TYPE (2              ),
   .S02_AW_REG_TYPE(0              ),
   .S02_W_REG_TYPE (0              ),
   .S02_B_REG_TYPE (1              ),
   .S02_AR_REG_TYPE(0              ),
   .S02_R_REG_TYPE (2              ),
   .M00_AW_REG_TYPE(1              ),
   .M00_W_REG_TYPE (2              ),
   .M00_B_REG_TYPE (0              ),
   .M00_AR_REG_TYPE(1              ),
   .M00_R_REG_TYPE (0              ),
   .M01_AW_REG_TYPE(1              ),
   .M01_W_REG_TYPE (2              ),
   .M01_B_REG_TYPE (0              ),
   .M01_AR_REG_TYPE(1              ),
   .M01_R_REG_TYPE (0              ),
   .M02_AW_REG_TYPE(1              ),
   .M02_W_REG_TYPE (2              ),
   .M02_B_REG_TYPE (0              ),
   .M02_AR_REG_TYPE(1              ),
   .M02_R_REG_TYPE (0              ),
   .M03_AW_REG_TYPE(1              ),
   .M03_W_REG_TYPE (2              ),
   .M03_B_REG_TYPE (0              ),
   .M03_AR_REG_TYPE(1              ),
   .M03_R_REG_TYPE (0              )
)
 u_axi_tmr_voter_ds_1m3s_inst1(
    .clk                                (clk                       ),
    .rst                                (rst                       ),
//s00
    .s00_axi_awid                       (s00_vd1_axi_awid              ),
    .s00_axi_awaddr                     (s00_vd1_axi_awaddr            ),
    .s00_axi_awlen                      (s00_vd1_axi_awlen             ),
    .s00_axi_awsize                     (s00_vd1_axi_awsize            ),
    .s00_axi_awburst                    (s00_vd1_axi_awburst           ),
    .s00_axi_awlock                     (s00_vd1_axi_awlock            ),
    .s00_axi_awcache                    (s00_vd1_axi_awcache           ),
    .s00_axi_awprot                     (s00_vd1_axi_awprot            ),
    .s00_axi_awqos                      (s00_vd1_axi_awqos             ),
    .s00_axi_awregion                   (s00_vd1_axi_awregion          ),
    .s00_axi_awuser                     (s00_vd1_axi_awuser            ),
    .s00_axi_awvalid                    (s00_vd1_axi_awvalid           ),
    .s00_axi_awready                    (s00_vd1_axi_awready           ),
    .s00_axi_wdata                      (s00_vd1_axi_wdata             ),
    .s00_axi_wstrb                      (s00_vd1_axi_wstrb             ),
    .s00_axi_wlast                      (s00_vd1_axi_wlast             ),
    .s00_axi_wuser                      (s00_vd1_axi_wuser             ),
    .s00_axi_wvalid                     (s00_vd1_axi_wvalid            ),
    .s00_axi_wready                     (s00_vd1_axi_wready            ),
    .s00_axi_bid                        (s00_vd1_axi_bid               ),
    .s00_axi_bresp                      (s00_vd1_axi_bresp             ),
    .s00_axi_buser                      (s00_vd1_axi_buser             ),
    .s00_axi_bvalid                     (s00_vd1_axi_bvalid            ),
    .s00_axi_bready                     (s00_vd1_axi_bready            ),
    .s00_axi_arid                       (s00_vd1_axi_arid              ),
    .s00_axi_araddr                     (s00_vd1_axi_araddr            ),
    .s00_axi_arlen                      (s00_vd1_axi_arlen             ),
    .s00_axi_arsize                     (s00_vd1_axi_arsize            ),
    .s00_axi_arburst                    (s00_vd1_axi_arburst           ),
    .s00_axi_arlock                     (s00_vd1_axi_arlock            ),
    .s00_axi_arcache                    (s00_vd1_axi_arcache           ),
    .s00_axi_arprot                     (s00_vd1_axi_arprot            ),
    .s00_axi_arqos                      (s00_vd1_axi_arqos             ),
    .s00_axi_arregion                   (s00_vd1_axi_arregion          ),
    .s00_axi_aruser                     (s00_vd1_axi_aruser            ),
    .s00_axi_arvalid                    (s00_vd1_axi_arvalid           ),
    .s00_axi_arready                    (s00_vd1_axi_arready           ),
    .s00_axi_rid                        (s00_vd1_axi_rid               ),
    .s00_axi_rdata                      (s00_vd1_axi_rdata             ),
    .s00_axi_rresp                      (s00_vd1_axi_rresp             ),
    .s00_axi_rlast                      (s00_vd1_axi_rlast             ),
    .s00_axi_ruser                      (s00_vd1_axi_ruser             ),
    .s00_axi_rvalid                     (s00_vd1_axi_rvalid            ),
    .s00_axi_rready                     (s00_vd1_axi_rready            ),
//s01
    .s01_axi_awid                       (s01_vd1_axi_awid              ),
    .s01_axi_awaddr                     (s01_vd1_axi_awaddr            ),
    .s01_axi_awlen                      (s01_vd1_axi_awlen             ),
    .s01_axi_awsize                     (s01_vd1_axi_awsize            ),
    .s01_axi_awburst                    (s01_vd1_axi_awburst           ),
    .s01_axi_awlock                     (s01_vd1_axi_awlock            ),
    .s01_axi_awcache                    (s01_vd1_axi_awcache           ),
    .s01_axi_awprot                     (s01_vd1_axi_awprot            ),
    .s01_axi_awqos                      (s01_vd1_axi_awqos             ),
    .s01_axi_awregion                   (s01_vd1_axi_awregion          ),
    .s01_axi_awuser                     (s01_vd1_axi_awuser            ),
    .s01_axi_awvalid                    (s01_vd1_axi_awvalid           ),
    .s01_axi_awready                    (s01_vd1_axi_awready           ),
    .s01_axi_wdata                      (s01_vd1_axi_wdata             ),
    .s01_axi_wstrb                      (s01_vd1_axi_wstrb             ),
    .s01_axi_wlast                      (s01_vd1_axi_wlast             ),
    .s01_axi_wuser                      (s01_vd1_axi_wuser             ),
    .s01_axi_wvalid                     (s01_vd1_axi_wvalid            ),
    .s01_axi_wready                     (s01_vd1_axi_wready            ),
    .s01_axi_bid                        (s01_vd1_axi_bid               ),
    .s01_axi_bresp                      (s01_vd1_axi_bresp             ),
    .s01_axi_buser                      (s01_vd1_axi_buser             ),
    .s01_axi_bvalid                     (s01_vd1_axi_bvalid            ),
    .s01_axi_bready                     (s01_vd1_axi_bready            ),
    .s01_axi_arid                       (s01_vd1_axi_arid              ),
    .s01_axi_araddr                     (s01_vd1_axi_araddr            ),
    .s01_axi_arlen                      (s01_vd1_axi_arlen             ),
    .s01_axi_arsize                     (s01_vd1_axi_arsize            ),
    .s01_axi_arburst                    (s01_vd1_axi_arburst           ),
    .s01_axi_arlock                     (s01_vd1_axi_arlock            ),
    .s01_axi_arcache                    (s01_vd1_axi_arcache           ),
    .s01_axi_arprot                     (s01_vd1_axi_arprot            ),
    .s01_axi_arqos                      (s01_vd1_axi_arqos             ),
    .s01_axi_arregion                   (s01_vd1_axi_arregion          ),
    .s01_axi_aruser                     (s01_vd1_axi_aruser            ),
    .s01_axi_arvalid                    (s01_vd1_axi_arvalid           ),
    .s01_axi_arready                    (s01_vd1_axi_arready           ),
    .s01_axi_rid                        (s01_vd1_axi_rid               ),
    .s01_axi_rdata                      (s01_vd1_axi_rdata             ),
    .s01_axi_rresp                      (s01_vd1_axi_rresp             ),
    .s01_axi_rlast                      (s01_vd1_axi_rlast             ),
    .s01_axi_ruser                      (s01_vd1_axi_ruser             ),
    .s01_axi_rvalid                     (s01_vd1_axi_rvalid            ),
    .s01_axi_rready                     (s01_vd1_axi_rready            ),
//s02
    .s02_axi_awid                       (s02_vd1_axi_awid              ),
    .s02_axi_awaddr                     (s02_vd1_axi_awaddr            ),
    .s02_axi_awlen                      (s02_vd1_axi_awlen             ),
    .s02_axi_awsize                     (s02_vd1_axi_awsize            ),
    .s02_axi_awburst                    (s02_vd1_axi_awburst           ),
    .s02_axi_awlock                     (s02_vd1_axi_awlock            ),
    .s02_axi_awcache                    (s02_vd1_axi_awcache           ),
    .s02_axi_awprot                     (s02_vd1_axi_awprot            ),
    .s02_axi_awqos                      (s02_vd1_axi_awqos             ),
    .s02_axi_awregion                   (s02_vd1_axi_awregion          ),
    .s02_axi_awuser                     (s02_vd1_axi_awuser            ),
    .s02_axi_awvalid                    (s02_vd1_axi_awvalid           ),
    .s02_axi_awready                    (s02_vd1_axi_awready           ),
    .s02_axi_wdata                      (s02_vd1_axi_wdata             ),
    .s02_axi_wstrb                      (s02_vd1_axi_wstrb             ),
    .s02_axi_wlast                      (s02_vd1_axi_wlast             ),
    .s02_axi_wuser                      (s02_vd1_axi_wuser             ),
    .s02_axi_wvalid                     (s02_vd1_axi_wvalid            ),
    .s02_axi_wready                     (s02_vd1_axi_wready            ),
    .s02_axi_bid                        (s02_vd1_axi_bid               ),
    .s02_axi_bresp                      (s02_vd1_axi_bresp             ),
    .s02_axi_buser                      (s02_vd1_axi_buser             ),
    .s02_axi_bvalid                     (s02_vd1_axi_bvalid            ),
    .s02_axi_bready                     (s02_vd1_axi_bready            ),
    .s02_axi_arid                       (s02_vd1_axi_arid              ),
    .s02_axi_araddr                     (s02_vd1_axi_araddr            ),
    .s02_axi_arlen                      (s02_vd1_axi_arlen             ),
    .s02_axi_arsize                     (s02_vd1_axi_arsize            ),
    .s02_axi_arburst                    (s02_vd1_axi_arburst           ),
    .s02_axi_arlock                     (s02_vd1_axi_arlock            ),
    .s02_axi_arcache                    (s02_vd1_axi_arcache           ),
    .s02_axi_arprot                     (s02_vd1_axi_arprot            ),
    .s02_axi_arqos                      (s02_vd1_axi_arqos             ),
    .s02_axi_arregion                   (s02_vd1_axi_arregion          ),
    .s02_axi_aruser                     (s02_vd1_axi_aruser            ),
    .s02_axi_arvalid                    (s02_vd1_axi_arvalid           ),
    .s02_axi_arready                    (s02_vd1_axi_arready           ),
    .s02_axi_rid                        (s02_vd1_axi_rid               ),
    .s02_axi_rdata                      (s02_vd1_axi_rdata             ),
    .s02_axi_rresp                      (s02_vd1_axi_rresp             ),
    .s02_axi_rlast                      (s02_vd1_axi_rlast             ),
    .s02_axi_ruser                      (s02_vd1_axi_ruser             ),
    .s02_axi_rvalid                     (s02_vd1_axi_rvalid            ),
    .s02_axi_rready                     (s02_vd1_axi_rready            ),
//m01
    .m00_axi_awid                       (m01_axi_awid              ),
    .m00_axi_awaddr                     (m01_axi_awaddr            ),
    .m00_axi_awlen                      (m01_axi_awlen             ),
    .m00_axi_awsize                     (m01_axi_awsize            ),
    .m00_axi_awburst                    (m01_axi_awburst           ),
    .m00_axi_awlock                     (m01_axi_awlock            ),
    .m00_axi_awcache                    (m01_axi_awcache           ),
    .m00_axi_awprot                     (m01_axi_awprot            ),
    .m00_axi_awqos                      (m01_axi_awqos             ),
    .m00_axi_awregion                   (m01_axi_awregion          ),
    .m00_axi_awuser                     (m01_axi_awuser            ),
    .m00_axi_awvalid                    (m01_axi_awvalid           ),
    .m00_axi_awready                    (m01_axi_awready           ),
    .m00_axi_wdata                      (m01_axi_wdata             ),
    .m00_axi_wstrb                      (m01_axi_wstrb             ),
    .m00_axi_wlast                      (m01_axi_wlast             ),
    .m00_axi_wuser                      (m01_axi_wuser             ),
    .m00_axi_wvalid                     (m01_axi_wvalid            ),
    .m00_axi_wready                     (m01_axi_wready            ),
    .m00_axi_bid                        (m01_axi_bid               ),
    .m00_axi_bresp                      (m01_axi_bresp             ),
    .m00_axi_buser                      (m01_axi_buser             ),
    .m00_axi_bvalid                     (m01_axi_bvalid            ),
    .m00_axi_bready                     (m01_axi_bready            ),
    .m00_axi_arid                       (m01_axi_arid              ),
    .m00_axi_araddr                     (m01_axi_araddr            ),
    .m00_axi_arlen                      (m01_axi_arlen             ),
    .m00_axi_arsize                     (m01_axi_arsize            ),
    .m00_axi_arburst                    (m01_axi_arburst           ),
    .m00_axi_arlock                     (m01_axi_arlock            ),
    .m00_axi_arcache                    (m01_axi_arcache           ),
    .m00_axi_arprot                     (m01_axi_arprot            ),
    .m00_axi_arqos                      (m01_axi_arqos             ),
    .m00_axi_arregion                   (m01_axi_arregion          ),
    .m00_axi_aruser                     (m01_axi_aruser            ),
    .m00_axi_arvalid                    (m01_axi_arvalid           ),
    .m00_axi_arready                    (m01_axi_arready           ),
    .m00_axi_rid                        (m01_axi_rid               ),
    .m00_axi_rdata                      (m01_axi_rdata             ),
    .m00_axi_rresp                      (m01_axi_rresp             ),
    .m00_axi_rlast                      (m01_axi_rlast             ),
    .m00_axi_ruser                      (m01_axi_ruser             ),
    .m00_axi_rvalid                     (m01_axi_rvalid            ),
    .m00_axi_rready                     (m01_axi_rready            )
);

//inst2
//m02+vd2
axi_tmr_voter_ds_1m3s#(
   .DATA_WIDTH     (64             ),
   .ADDR_WIDTH     (32             ),
   .STRB_WIDTH     ((DATA_WIDTH/8) ),
   .S_ID_WIDTH     (8              ),
   .M_ID_WIDTH     (S_ID_WIDTH+$clog2(3)),
   .AWUSER_ENABLE  (0              ),
   .AWUSER_WIDTH   (1              ),
   .WUSER_ENABLE   (0              ),
   .WUSER_WIDTH    (1              ),
   .BUSER_ENABLE   (0              ),
   .BUSER_WIDTH    (1              ),
   .ARUSER_ENABLE  (0              ),
   .ARUSER_WIDTH   (1              ),
   .RUSER_ENABLE   (0              ),
   .RUSER_WIDTH    (1              ),
   .S00_THREADS    (8              ),
   .S00_ACCEPT     (16             ),
   .S01_THREADS    (8              ),
   .S01_ACCEPT     (16             ),
   .S02_THREADS    (8              ),
   .S02_ACCEPT     (16             ),
   .M_REGIONS      (1              ),
   .M00_BASE_ADDR  (0              ),
   .M00_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M00_CONNECT_READ(3'b100         ),
   .M00_CONNECT_WRITE(3'b100         ),
   .M00_ISSUE      (8              ),
   .M00_SECURE     (1              ),
   .M01_BASE_ADDR  (0              ),
   .M01_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M01_CONNECT_READ(3'b011         ),
   .M01_CONNECT_WRITE(3'b011         ),
   .M01_ISSUE      (8              ),
   .M01_SECURE     (0              ),
   .M02_BASE_ADDR  (0              ),
   .M02_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M02_CONNECT_READ(3'b100         ),
   .M02_CONNECT_WRITE(3'b100         ),
   .M02_ISSUE      (8              ),
   .M02_SECURE     (1              ),
   .M03_BASE_ADDR  (0              ),
   .M03_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M03_CONNECT_READ(3'b011         ),
   .M03_CONNECT_WRITE(3'b011         ),
   .M03_ISSUE      (8              ),
   .M03_SECURE     (0              ),
   .S00_AW_REG_TYPE(0              ),
   .S00_W_REG_TYPE (0              ),
   .S00_B_REG_TYPE (1              ),
   .S00_AR_REG_TYPE(0              ),
   .S00_R_REG_TYPE (2              ),
   .S01_AW_REG_TYPE(0              ),
   .S01_W_REG_TYPE (0              ),
   .S01_B_REG_TYPE (1              ),
   .S01_AR_REG_TYPE(0              ),
   .S01_R_REG_TYPE (2              ),
   .S02_AW_REG_TYPE(0              ),
   .S02_W_REG_TYPE (0              ),
   .S02_B_REG_TYPE (1              ),
   .S02_AR_REG_TYPE(0              ),
   .S02_R_REG_TYPE (2              ),
   .M00_AW_REG_TYPE(1              ),
   .M00_W_REG_TYPE (2              ),
   .M00_B_REG_TYPE (0              ),
   .M00_AR_REG_TYPE(1              ),
   .M00_R_REG_TYPE (0              ),
   .M01_AW_REG_TYPE(1              ),
   .M01_W_REG_TYPE (2              ),
   .M01_B_REG_TYPE (0              ),
   .M01_AR_REG_TYPE(1              ),
   .M01_R_REG_TYPE (0              ),
   .M02_AW_REG_TYPE(1              ),
   .M02_W_REG_TYPE (2              ),
   .M02_B_REG_TYPE (0              ),
   .M02_AR_REG_TYPE(1              ),
   .M02_R_REG_TYPE (0              ),
   .M03_AW_REG_TYPE(1              ),
   .M03_W_REG_TYPE (2              ),
   .M03_B_REG_TYPE (0              ),
   .M03_AR_REG_TYPE(1              ),
   .M03_R_REG_TYPE (0              )
)
 u_axi_tmr_voter_ds_1m3s_inst2(
    .clk                                (clk                       ),
    .rst                                (rst                       ),
//s00
    .s00_axi_awid                       (s00_vd2_axi_awid              ),
    .s00_axi_awaddr                     (s00_vd2_axi_awaddr            ),
    .s00_axi_awlen                      (s00_vd2_axi_awlen             ),
    .s00_axi_awsize                     (s00_vd2_axi_awsize            ),
    .s00_axi_awburst                    (s00_vd2_axi_awburst           ),
    .s00_axi_awlock                     (s00_vd2_axi_awlock            ),
    .s00_axi_awcache                    (s00_vd2_axi_awcache           ),
    .s00_axi_awprot                     (s00_vd2_axi_awprot            ),
    .s00_axi_awqos                      (s00_vd2_axi_awqos             ),
    .s00_axi_awregion                   (s00_vd2_axi_awregion          ),
    .s00_axi_awuser                     (s00_vd2_axi_awuser            ),
    .s00_axi_awvalid                    (s00_vd2_axi_awvalid           ),
    .s00_axi_awready                    (s00_vd2_axi_awready           ),
    .s00_axi_wdata                      (s00_vd2_axi_wdata             ),
    .s00_axi_wstrb                      (s00_vd2_axi_wstrb             ),
    .s00_axi_wlast                      (s00_vd2_axi_wlast             ),
    .s00_axi_wuser                      (s00_vd2_axi_wuser             ),
    .s00_axi_wvalid                     (s00_vd2_axi_wvalid            ),
    .s00_axi_wready                     (s00_vd2_axi_wready            ),
    .s00_axi_bid                        (s00_vd2_axi_bid               ),
    .s00_axi_bresp                      (s00_vd2_axi_bresp             ),
    .s00_axi_buser                      (s00_vd2_axi_buser             ),
    .s00_axi_bvalid                     (s00_vd2_axi_bvalid            ),
    .s00_axi_bready                     (s00_vd2_axi_bready            ),
    .s00_axi_arid                       (s00_vd2_axi_arid              ),
    .s00_axi_araddr                     (s00_vd2_axi_araddr            ),
    .s00_axi_arlen                      (s00_vd2_axi_arlen             ),
    .s00_axi_arsize                     (s00_vd2_axi_arsize            ),
    .s00_axi_arburst                    (s00_vd2_axi_arburst           ),
    .s00_axi_arlock                     (s00_vd2_axi_arlock            ),
    .s00_axi_arcache                    (s00_vd2_axi_arcache           ),
    .s00_axi_arprot                     (s00_vd2_axi_arprot            ),
    .s00_axi_arqos                      (s00_vd2_axi_arqos             ),
    .s00_axi_arregion                   (s00_vd2_axi_arregion          ),
    .s00_axi_aruser                     (s00_vd2_axi_aruser            ),
    .s00_axi_arvalid                    (s00_vd2_axi_arvalid           ),
    .s00_axi_arready                    (s00_vd2_axi_arready           ),
    .s00_axi_rid                        (s00_vd2_axi_rid               ),
    .s00_axi_rdata                      (s00_vd2_axi_rdata             ),
    .s00_axi_rresp                      (s00_vd2_axi_rresp             ),
    .s00_axi_rlast                      (s00_vd2_axi_rlast             ),
    .s00_axi_ruser                      (s00_vd2_axi_ruser             ),
    .s00_axi_rvalid                     (s00_vd2_axi_rvalid            ),
    .s00_axi_rready                     (s00_vd2_axi_rready            ),
//s01
    .s01_axi_awid                       (s01_vd2_axi_awid              ),
    .s01_axi_awaddr                     (s01_vd2_axi_awaddr            ),
    .s01_axi_awlen                      (s01_vd2_axi_awlen             ),
    .s01_axi_awsize                     (s01_vd2_axi_awsize            ),
    .s01_axi_awburst                    (s01_vd2_axi_awburst           ),
    .s01_axi_awlock                     (s01_vd2_axi_awlock            ),
    .s01_axi_awcache                    (s01_vd2_axi_awcache           ),
    .s01_axi_awprot                     (s01_vd2_axi_awprot            ),
    .s01_axi_awqos                      (s01_vd2_axi_awqos             ),
    .s01_axi_awregion                   (s01_vd2_axi_awregion          ),
    .s01_axi_awuser                     (s01_vd2_axi_awuser            ),
    .s01_axi_awvalid                    (s01_vd2_axi_awvalid           ),
    .s01_axi_awready                    (s01_vd2_axi_awready           ),
    .s01_axi_wdata                      (s01_vd2_axi_wdata             ),
    .s01_axi_wstrb                      (s01_vd2_axi_wstrb             ),
    .s01_axi_wlast                      (s01_vd2_axi_wlast             ),
    .s01_axi_wuser                      (s01_vd2_axi_wuser             ),
    .s01_axi_wvalid                     (s01_vd2_axi_wvalid            ),
    .s01_axi_wready                     (s01_vd2_axi_wready            ),
    .s01_axi_bid                        (s01_vd2_axi_bid               ),
    .s01_axi_bresp                      (s01_vd2_axi_bresp             ),
    .s01_axi_buser                      (s01_vd2_axi_buser             ),
    .s01_axi_bvalid                     (s01_vd2_axi_bvalid            ),
    .s01_axi_bready                     (s01_vd2_axi_bready            ),
    .s01_axi_arid                       (s01_vd2_axi_arid              ),
    .s01_axi_araddr                     (s01_vd2_axi_araddr            ),
    .s01_axi_arlen                      (s01_vd2_axi_arlen             ),
    .s01_axi_arsize                     (s01_vd2_axi_arsize            ),
    .s01_axi_arburst                    (s01_vd2_axi_arburst           ),
    .s01_axi_arlock                     (s01_vd2_axi_arlock            ),
    .s01_axi_arcache                    (s01_vd2_axi_arcache           ),
    .s01_axi_arprot                     (s01_vd2_axi_arprot            ),
    .s01_axi_arqos                      (s01_vd2_axi_arqos             ),
    .s01_axi_arregion                   (s01_vd2_axi_arregion          ),
    .s01_axi_aruser                     (s01_vd2_axi_aruser            ),
    .s01_axi_arvalid                    (s01_vd2_axi_arvalid           ),
    .s01_axi_arready                    (s01_vd2_axi_arready           ),
    .s01_axi_rid                        (s01_vd2_axi_rid               ),
    .s01_axi_rdata                      (s01_vd2_axi_rdata             ),
    .s01_axi_rresp                      (s01_vd2_axi_rresp             ),
    .s01_axi_rlast                      (s01_vd2_axi_rlast             ),
    .s01_axi_ruser                      (s01_vd2_axi_ruser             ),
    .s01_axi_rvalid                     (s01_vd2_axi_rvalid            ),
    .s01_axi_rready                     (s01_vd2_axi_rready            ),
//s02
    .s02_axi_awid                       (s02_vd2_axi_awid              ),
    .s02_axi_awaddr                     (s02_vd2_axi_awaddr            ),
    .s02_axi_awlen                      (s02_vd2_axi_awlen             ),
    .s02_axi_awsize                     (s02_vd2_axi_awsize            ),
    .s02_axi_awburst                    (s02_vd2_axi_awburst           ),
    .s02_axi_awlock                     (s02_vd2_axi_awlock            ),
    .s02_axi_awcache                    (s02_vd2_axi_awcache           ),
    .s02_axi_awprot                     (s02_vd2_axi_awprot            ),
    .s02_axi_awqos                      (s02_vd2_axi_awqos             ),
    .s02_axi_awregion                   (s02_vd2_axi_awregion          ),
    .s02_axi_awuser                     (s02_vd2_axi_awuser            ),
    .s02_axi_awvalid                    (s02_vd2_axi_awvalid           ),
    .s02_axi_awready                    (s02_vd2_axi_awready           ),
    .s02_axi_wdata                      (s02_vd2_axi_wdata             ),
    .s02_axi_wstrb                      (s02_vd2_axi_wstrb             ),
    .s02_axi_wlast                      (s02_vd2_axi_wlast             ),
    .s02_axi_wuser                      (s02_vd2_axi_wuser             ),
    .s02_axi_wvalid                     (s02_vd2_axi_wvalid            ),
    .s02_axi_wready                     (s02_vd2_axi_wready            ),
    .s02_axi_bid                        (s02_vd2_axi_bid               ),
    .s02_axi_bresp                      (s02_vd2_axi_bresp             ),
    .s02_axi_buser                      (s02_vd2_axi_buser             ),
    .s02_axi_bvalid                     (s02_vd2_axi_bvalid            ),
    .s02_axi_bready                     (s02_vd2_axi_bready            ),
    .s02_axi_arid                       (s02_vd2_axi_arid              ),
    .s02_axi_araddr                     (s02_vd2_axi_araddr            ),
    .s02_axi_arlen                      (s02_vd2_axi_arlen             ),
    .s02_axi_arsize                     (s02_vd2_axi_arsize            ),
    .s02_axi_arburst                    (s02_vd2_axi_arburst           ),
    .s02_axi_arlock                     (s02_vd2_axi_arlock            ),
    .s02_axi_arcache                    (s02_vd2_axi_arcache           ),
    .s02_axi_arprot                     (s02_vd2_axi_arprot            ),
    .s02_axi_arqos                      (s02_vd2_axi_arqos             ),
    .s02_axi_arregion                   (s02_vd2_axi_arregion          ),
    .s02_axi_aruser                     (s02_vd2_axi_aruser            ),
    .s02_axi_arvalid                    (s02_vd2_axi_arvalid           ),
    .s02_axi_arready                    (s02_vd2_axi_arready           ),
    .s02_axi_rid                        (s02_vd2_axi_rid               ),
    .s02_axi_rdata                      (s02_vd2_axi_rdata             ),
    .s02_axi_rresp                      (s02_vd2_axi_rresp             ),
    .s02_axi_rlast                      (s02_vd2_axi_rlast             ),
    .s02_axi_ruser                      (s02_vd2_axi_ruser             ),
    .s02_axi_rvalid                     (s02_vd2_axi_rvalid            ),
    .s02_axi_rready                     (s02_vd2_axi_rready            ),
//m02
    .m00_axi_awid                       (m02_axi_awid              ),
    .m00_axi_awaddr                     (m02_axi_awaddr            ),
    .m00_axi_awlen                      (m02_axi_awlen             ),
    .m00_axi_awsize                     (m02_axi_awsize            ),
    .m00_axi_awburst                    (m02_axi_awburst           ),
    .m00_axi_awlock                     (m02_axi_awlock            ),
    .m00_axi_awcache                    (m02_axi_awcache           ),
    .m00_axi_awprot                     (m02_axi_awprot            ),
    .m00_axi_awqos                      (m02_axi_awqos             ),
    .m00_axi_awregion                   (m02_axi_awregion          ),
    .m00_axi_awuser                     (m02_axi_awuser            ),
    .m00_axi_awvalid                    (m02_axi_awvalid           ),
    .m00_axi_awready                    (m02_axi_awready           ),
    .m00_axi_wdata                      (m02_axi_wdata             ),
    .m00_axi_wstrb                      (m02_axi_wstrb             ),
    .m00_axi_wlast                      (m02_axi_wlast             ),
    .m00_axi_wuser                      (m02_axi_wuser             ),
    .m00_axi_wvalid                     (m02_axi_wvalid            ),
    .m00_axi_wready                     (m02_axi_wready            ),
    .m00_axi_bid                        (m02_axi_bid               ),
    .m00_axi_bresp                      (m02_axi_bresp             ),
    .m00_axi_buser                      (m02_axi_buser             ),
    .m00_axi_bvalid                     (m02_axi_bvalid            ),
    .m00_axi_bready                     (m02_axi_bready            ),
    .m00_axi_arid                       (m02_axi_arid              ),
    .m00_axi_araddr                     (m02_axi_araddr            ),
    .m00_axi_arlen                      (m02_axi_arlen             ),
    .m00_axi_arsize                     (m02_axi_arsize            ),
    .m00_axi_arburst                    (m02_axi_arburst           ),
    .m00_axi_arlock                     (m02_axi_arlock            ),
    .m00_axi_arcache                    (m02_axi_arcache           ),
    .m00_axi_arprot                     (m02_axi_arprot            ),
    .m00_axi_arqos                      (m02_axi_arqos             ),
    .m00_axi_arregion                   (m02_axi_arregion          ),
    .m00_axi_aruser                     (m02_axi_aruser            ),
    .m00_axi_arvalid                    (m02_axi_arvalid           ),
    .m00_axi_arready                    (m02_axi_arready           ),
    .m00_axi_rid                        (m02_axi_rid               ),
    .m00_axi_rdata                      (m02_axi_rdata             ),
    .m00_axi_rresp                      (m02_axi_rresp             ),
    .m00_axi_rlast                      (m02_axi_rlast             ),
    .m00_axi_ruser                      (m02_axi_ruser             ),
    .m00_axi_rvalid                     (m02_axi_rvalid            ),
    .m00_axi_rready                     (m02_axi_rready            )
);

//inst3
//m03+vd3
axi_tmr_voter_ds_1m3s#(
   .DATA_WIDTH     (64             ),
   .ADDR_WIDTH     (32             ),
   .STRB_WIDTH     ((DATA_WIDTH/8) ),
   .S_ID_WIDTH     (8              ),
   .M_ID_WIDTH     (S_ID_WIDTH+$clog2(3)),
   .AWUSER_ENABLE  (0              ),
   .AWUSER_WIDTH   (1              ),
   .WUSER_ENABLE   (0              ),
   .WUSER_WIDTH    (1              ),
   .BUSER_ENABLE   (0              ),
   .BUSER_WIDTH    (1              ),
   .ARUSER_ENABLE  (0              ),
   .ARUSER_WIDTH   (1              ),
   .RUSER_ENABLE   (0              ),
   .RUSER_WIDTH    (1              ),
   .S00_THREADS    (8              ),
   .S00_ACCEPT     (16             ),
   .S01_THREADS    (8              ),
   .S01_ACCEPT     (16             ),
   .S02_THREADS    (8              ),
   .S02_ACCEPT     (16             ),
   .M_REGIONS      (1              ),
   .M00_BASE_ADDR  (0              ),
   .M00_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M00_CONNECT_READ(3'b100         ),
   .M00_CONNECT_WRITE(3'b100         ),
   .M00_ISSUE      (8              ),
   .M00_SECURE     (1              ),
   .M01_BASE_ADDR  (0              ),
   .M01_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M01_CONNECT_READ(3'b011         ),
   .M01_CONNECT_WRITE(3'b011         ),
   .M01_ISSUE      (8              ),
   .M01_SECURE     (0              ),
   .M02_BASE_ADDR  (0              ),
   .M02_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M02_CONNECT_READ(3'b100         ),
   .M02_CONNECT_WRITE(3'b100         ),
   .M02_ISSUE      (8              ),
   .M02_SECURE     (1              ),
   .M03_BASE_ADDR  (0              ),
   .M03_ADDR_WIDTH ({M_REGIONS{32'd24}}),
   .M03_CONNECT_READ(3'b011         ),
   .M03_CONNECT_WRITE(3'b011         ),
   .M03_ISSUE      (8              ),
   .M03_SECURE     (0              ),
   .S00_AW_REG_TYPE(0              ),
   .S00_W_REG_TYPE (0              ),
   .S00_B_REG_TYPE (1              ),
   .S00_AR_REG_TYPE(0              ),
   .S00_R_REG_TYPE (2              ),
   .S01_AW_REG_TYPE(0              ),
   .S01_W_REG_TYPE (0              ),
   .S01_B_REG_TYPE (1              ),
   .S01_AR_REG_TYPE(0              ),
   .S01_R_REG_TYPE (2              ),
   .S02_AW_REG_TYPE(0              ),
   .S02_W_REG_TYPE (0              ),
   .S02_B_REG_TYPE (1              ),
   .S02_AR_REG_TYPE(0              ),
   .S02_R_REG_TYPE (2              ),
   .M00_AW_REG_TYPE(1              ),
   .M00_W_REG_TYPE (2              ),
   .M00_B_REG_TYPE (0              ),
   .M00_AR_REG_TYPE(1              ),
   .M00_R_REG_TYPE (0              ),
   .M01_AW_REG_TYPE(1              ),
   .M01_W_REG_TYPE (2              ),
   .M01_B_REG_TYPE (0              ),
   .M01_AR_REG_TYPE(1              ),
   .M01_R_REG_TYPE (0              ),
   .M02_AW_REG_TYPE(1              ),
   .M02_W_REG_TYPE (2              ),
   .M02_B_REG_TYPE (0              ),
   .M02_AR_REG_TYPE(1              ),
   .M02_R_REG_TYPE (0              ),
   .M03_AW_REG_TYPE(1              ),
   .M03_W_REG_TYPE (2              ),
   .M03_B_REG_TYPE (0              ),
   .M03_AR_REG_TYPE(1              ),
   .M03_R_REG_TYPE (0              )
)
 u_axi_tmr_voter_ds_1m3s_inst3(
    .clk                                (clk                       ),
    .rst                                (rst                       ),
//s00
    .s00_axi_awid                       (s00_vd3_axi_awid              ),
    .s00_axi_awaddr                     (s00_vd3_axi_awaddr            ),
    .s00_axi_awlen                      (s00_vd3_axi_awlen             ),
    .s00_axi_awsize                     (s00_vd3_axi_awsize            ),
    .s00_axi_awburst                    (s00_vd3_axi_awburst           ),
    .s00_axi_awlock                     (s00_vd3_axi_awlock            ),
    .s00_axi_awcache                    (s00_vd3_axi_awcache           ),
    .s00_axi_awprot                     (s00_vd3_axi_awprot            ),
    .s00_axi_awqos                      (s00_vd3_axi_awqos             ),
    .s00_axi_awregion                   (s00_vd3_axi_awregion          ),
    .s00_axi_awuser                     (s00_vd3_axi_awuser            ),
    .s00_axi_awvalid                    (s00_vd3_axi_awvalid           ),
    .s00_axi_awready                    (s00_vd3_axi_awready           ),
    .s00_axi_wdata                      (s00_vd3_axi_wdata             ),
    .s00_axi_wstrb                      (s00_vd3_axi_wstrb             ),
    .s00_axi_wlast                      (s00_vd3_axi_wlast             ),
    .s00_axi_wuser                      (s00_vd3_axi_wuser             ),
    .s00_axi_wvalid                     (s00_vd3_axi_wvalid            ),
    .s00_axi_wready                     (s00_vd3_axi_wready            ),
    .s00_axi_bid                        (s00_vd3_axi_bid               ),
    .s00_axi_bresp                      (s00_vd3_axi_bresp             ),
    .s00_axi_buser                      (s00_vd3_axi_buser             ),
    .s00_axi_bvalid                     (s00_vd3_axi_bvalid            ),
    .s00_axi_bready                     (s00_vd3_axi_bready            ),
    .s00_axi_arid                       (s00_vd3_axi_arid              ),
    .s00_axi_araddr                     (s00_vd3_axi_araddr            ),
    .s00_axi_arlen                      (s00_vd3_axi_arlen             ),
    .s00_axi_arsize                     (s00_vd3_axi_arsize            ),
    .s00_axi_arburst                    (s00_vd3_axi_arburst           ),
    .s00_axi_arlock                     (s00_vd3_axi_arlock            ),
    .s00_axi_arcache                    (s00_vd3_axi_arcache           ),
    .s00_axi_arprot                     (s00_vd3_axi_arprot            ),
    .s00_axi_arqos                      (s00_vd3_axi_arqos             ),
    .s00_axi_arregion                   (s00_vd3_axi_arregion          ),
    .s00_axi_aruser                     (s00_vd3_axi_aruser            ),
    .s00_axi_arvalid                    (s00_vd3_axi_arvalid           ),
    .s00_axi_arready                    (s00_vd3_axi_arready           ),
    .s00_axi_rid                        (s00_vd3_axi_rid               ),
    .s00_axi_rdata                      (s00_vd3_axi_rdata             ),
    .s00_axi_rresp                      (s00_vd3_axi_rresp             ),
    .s00_axi_rlast                      (s00_vd3_axi_rlast             ),
    .s00_axi_ruser                      (s00_vd3_axi_ruser             ),
    .s00_axi_rvalid                     (s00_vd3_axi_rvalid            ),
    .s00_axi_rready                     (s00_vd3_axi_rready            ),
//s01
    .s01_axi_awid                       (s01_vd3_axi_awid              ),
    .s01_axi_awaddr                     (s01_vd3_axi_awaddr            ),
    .s01_axi_awlen                      (s01_vd3_axi_awlen             ),
    .s01_axi_awsize                     (s01_vd3_axi_awsize            ),
    .s01_axi_awburst                    (s01_vd3_axi_awburst           ),
    .s01_axi_awlock                     (s01_vd3_axi_awlock            ),
    .s01_axi_awcache                    (s01_vd3_axi_awcache           ),
    .s01_axi_awprot                     (s01_vd3_axi_awprot            ),
    .s01_axi_awqos                      (s01_vd3_axi_awqos             ),
    .s01_axi_awregion                   (s01_vd3_axi_awregion          ),
    .s01_axi_awuser                     (s01_vd3_axi_awuser            ),
    .s01_axi_awvalid                    (s01_vd3_axi_awvalid           ),
    .s01_axi_awready                    (s01_vd3_axi_awready           ),
    .s01_axi_wdata                      (s01_vd3_axi_wdata             ),
    .s01_axi_wstrb                      (s01_vd3_axi_wstrb             ),
    .s01_axi_wlast                      (s01_vd3_axi_wlast             ),
    .s01_axi_wuser                      (s01_vd3_axi_wuser             ),
    .s01_axi_wvalid                     (s01_vd3_axi_wvalid            ),
    .s01_axi_wready                     (s01_vd3_axi_wready            ),
    .s01_axi_bid                        (s01_vd3_axi_bid               ),
    .s01_axi_bresp                      (s01_vd3_axi_bresp             ),
    .s01_axi_buser                      (s01_vd3_axi_buser             ),
    .s01_axi_bvalid                     (s01_vd3_axi_bvalid            ),
    .s01_axi_bready                     (s01_vd3_axi_bready            ),
    .s01_axi_arid                       (s01_vd3_axi_arid              ),
    .s01_axi_araddr                     (s01_vd3_axi_araddr            ),
    .s01_axi_arlen                      (s01_vd3_axi_arlen             ),
    .s01_axi_arsize                     (s01_vd3_axi_arsize            ),
    .s01_axi_arburst                    (s01_vd3_axi_arburst           ),
    .s01_axi_arlock                     (s01_vd3_axi_arlock            ),
    .s01_axi_arcache                    (s01_vd3_axi_arcache           ),
    .s01_axi_arprot                     (s01_vd3_axi_arprot            ),
    .s01_axi_arqos                      (s01_vd3_axi_arqos             ),
    .s01_axi_arregion                   (s01_vd3_axi_arregion          ),
    .s01_axi_aruser                     (s01_vd3_axi_aruser            ),
    .s01_axi_arvalid                    (s01_vd3_axi_arvalid           ),
    .s01_axi_arready                    (s01_vd3_axi_arready           ),
    .s01_axi_rid                        (s01_vd3_axi_rid               ),
    .s01_axi_rdata                      (s01_vd3_axi_rdata             ),
    .s01_axi_rresp                      (s01_vd3_axi_rresp             ),
    .s01_axi_rlast                      (s01_vd3_axi_rlast             ),
    .s01_axi_ruser                      (s01_vd3_axi_ruser             ),
    .s01_axi_rvalid                     (s01_vd3_axi_rvalid            ),
    .s01_axi_rready                     (s01_vd3_axi_rready            ),
//s02
    .s02_axi_awid                       (s02_vd3_axi_awid              ),
    .s02_axi_awaddr                     (s02_vd3_axi_awaddr            ),
    .s02_axi_awlen                      (s02_vd3_axi_awlen             ),
    .s02_axi_awsize                     (s02_vd3_axi_awsize            ),
    .s02_axi_awburst                    (s02_vd3_axi_awburst           ),
    .s02_axi_awlock                     (s02_vd3_axi_awlock            ),
    .s02_axi_awcache                    (s02_vd3_axi_awcache           ),
    .s02_axi_awprot                     (s02_vd3_axi_awprot            ),
    .s02_axi_awqos                      (s02_vd3_axi_awqos             ),
    .s02_axi_awregion                   (s02_vd3_axi_awregion          ),
    .s02_axi_awuser                     (s02_vd3_axi_awuser            ),
    .s02_axi_awvalid                    (s02_vd3_axi_awvalid           ),
    .s02_axi_awready                    (s02_vd3_axi_awready           ),
    .s02_axi_wdata                      (s02_vd3_axi_wdata             ),
    .s02_axi_wstrb                      (s02_vd3_axi_wstrb             ),
    .s02_axi_wlast                      (s02_vd3_axi_wlast             ),
    .s02_axi_wuser                      (s02_vd3_axi_wuser             ),
    .s02_axi_wvalid                     (s02_vd3_axi_wvalid            ),
    .s02_axi_wready                     (s02_vd3_axi_wready            ),
    .s02_axi_bid                        (s02_vd3_axi_bid               ),
    .s02_axi_bresp                      (s02_vd3_axi_bresp             ),
    .s02_axi_buser                      (s02_vd3_axi_buser             ),
    .s02_axi_bvalid                     (s02_vd3_axi_bvalid            ),
    .s02_axi_bready                     (s02_vd3_axi_bready            ),
    .s02_axi_arid                       (s02_vd3_axi_arid              ),
    .s02_axi_araddr                     (s02_vd3_axi_araddr            ),
    .s02_axi_arlen                      (s02_vd3_axi_arlen             ),
    .s02_axi_arsize                     (s02_vd3_axi_arsize            ),
    .s02_axi_arburst                    (s02_vd3_axi_arburst           ),
    .s02_axi_arlock                     (s02_vd3_axi_arlock            ),
    .s02_axi_arcache                    (s02_vd3_axi_arcache           ),
    .s02_axi_arprot                     (s02_vd3_axi_arprot            ),
    .s02_axi_arqos                      (s02_vd3_axi_arqos             ),
    .s02_axi_arregion                   (s02_vd3_axi_arregion          ),
    .s02_axi_aruser                     (s02_vd3_axi_aruser            ),
    .s02_axi_arvalid                    (s02_vd3_axi_arvalid           ),
    .s02_axi_arready                    (s02_vd3_axi_arready           ),
    .s02_axi_rid                        (s02_vd3_axi_rid               ),
    .s02_axi_rdata                      (s02_vd3_axi_rdata             ),
    .s02_axi_rresp                      (s02_vd3_axi_rresp             ),
    .s02_axi_rlast                      (s02_vd3_axi_rlast             ),
    .s02_axi_ruser                      (s02_vd3_axi_ruser             ),
    .s02_axi_rvalid                     (s02_vd3_axi_rvalid            ),
    .s02_axi_rready                     (s02_vd3_axi_rready            ),
//m03
    .m00_axi_awid                       (m03_axi_awid              ),
    .m00_axi_awaddr                     (m03_axi_awaddr            ),
    .m00_axi_awlen                      (m03_axi_awlen             ),
    .m00_axi_awsize                     (m03_axi_awsize            ),
    .m00_axi_awburst                    (m03_axi_awburst           ),
    .m00_axi_awlock                     (m03_axi_awlock            ),
    .m00_axi_awcache                    (m03_axi_awcache           ),
    .m00_axi_awprot                     (m03_axi_awprot            ),
    .m00_axi_awqos                      (m03_axi_awqos             ),
    .m00_axi_awregion                   (m03_axi_awregion          ),
    .m00_axi_awuser                     (m03_axi_awuser            ),
    .m00_axi_awvalid                    (m03_axi_awvalid           ),
    .m00_axi_awready                    (m03_axi_awready           ),
    .m00_axi_wdata                      (m03_axi_wdata             ),
    .m00_axi_wstrb                      (m03_axi_wstrb             ),
    .m00_axi_wlast                      (m03_axi_wlast             ),
    .m00_axi_wuser                      (m03_axi_wuser             ),
    .m00_axi_wvalid                     (m03_axi_wvalid            ),
    .m00_axi_wready                     (m03_axi_wready            ),
    .m00_axi_bid                        (m03_axi_bid               ),
    .m00_axi_bresp                      (m03_axi_bresp             ),
    .m00_axi_buser                      (m03_axi_buser             ),
    .m00_axi_bvalid                     (m03_axi_bvalid            ),
    .m00_axi_bready                     (m03_axi_bready            ),
    .m00_axi_arid                       (m03_axi_arid              ),
    .m00_axi_araddr                     (m03_axi_araddr            ),
    .m00_axi_arlen                      (m03_axi_arlen             ),
    .m00_axi_arsize                     (m03_axi_arsize            ),
    .m00_axi_arburst                    (m03_axi_arburst           ),
    .m00_axi_arlock                     (m03_axi_arlock            ),
    .m00_axi_arcache                    (m03_axi_arcache           ),
    .m00_axi_arprot                     (m03_axi_arprot            ),
    .m00_axi_arqos                      (m03_axi_arqos             ),
    .m00_axi_arregion                   (m03_axi_arregion          ),
    .m00_axi_aruser                     (m03_axi_aruser            ),
    .m00_axi_arvalid                    (m03_axi_arvalid           ),
    .m00_axi_arready                    (m03_axi_arready           ),
    .m00_axi_rid                        (m03_axi_rid               ),
    .m00_axi_rdata                      (m03_axi_rdata             ),
    .m00_axi_rresp                      (m03_axi_rresp             ),
    .m00_axi_rlast                      (m03_axi_rlast             ),
    .m00_axi_ruser                      (m03_axi_ruser             ),
    .m00_axi_rvalid                     (m03_axi_rvalid            ),
    .m00_axi_rready                     (m03_axi_rready            )
);
endmodule

`resetall
