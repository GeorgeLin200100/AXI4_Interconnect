`define AXI_AWID_IDX 1
`define AXI_AWADDR_IDX 2
`define AXI_AWLEN_IDX 3
`define AXI_AWSIZE_IDX 4
`define AXI_AWBURST_IDX 5
`define AXI_AWLOCK_IDX 6
`define AXI_AWCACHE_IDX 7
`define AXI_AWPROT_IDX 8
`define AXI_AWQOS_IDX 9
`define AXI_AWREGION_IDX 10
`define AXI_AWUSER_IDX 11
`define AXI_AWVALID_IDX 12
`define AXI_AWREADY_IDX 13
`define AXI_WDATA_IDX 14
`define AXI_WSTRB_IDX 15
`define AXI_WLAST_IDX 16
`define AXI_WUSER_IDX 17
`define AXI_WVALID_IDX 18
`define AXI_WREADY_IDX 19
`define AXI_BID_IDX 20
`define AXI_BRESP_IDX 21
`define AXI_BUSER_IDX 22
`define AXI_BVALID_IDX 23
`define AXI_BREADY_IDX 24
`define AXI_ARID_IDX 25
`define AXI_ARADDR_IDX 26
`define AXI_ARLEN_IDX 27
`define AXI_ARSIZE_IDX 28
`define AXI_ARBURST_IDX 29
`define AXI_ARLOCK_IDX 30
`define AXI_ARCACHE_IDX 31
`define AXI_ARPROT_IDX 32
`define AXI_ARQOS_IDX 33
`define AXI_ARREGION_IDX 34
`define AXI_ARUSER_IDX 35
`define AXI_ARVALID_IDX 36
`define AXI_ARREADY_IDX 37
`define AXI_RID_IDX 38
`define AXI_RDATA_IDX 39
`define AXI_RRESP_IDX 40
`define AXI_RLAST_IDX 41
`define AXI_RUSER_IDX 42
`define AXI_RVALID_IDX 43
`define AXI_RREADY_IDX 44