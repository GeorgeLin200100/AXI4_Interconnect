`ifndef TVIP_AXI_DEFINES_SVH
`define TVIP_AXI_DEFINES_SVH

`ifndef TVIP_AXI_MAX_ID_WIDTH
  //`define TVIP_AXI_MAX_ID_WIDTH 32
  define TVIP_AXI_MAX_ID_WIDTH 8
`endif

`ifndef TVIP_AXI_MAX_ADDRESS_WIDTH
  //`define TVIP_AXI_MAX_ADDRESS_WIDTH  64
  `define TVIP_AXI_MAX_ADDRESS_WIDTH  32
`endif

`ifndef TVIP_AXI_MAX_DATA_WIDTH
  //`define TVIP_AXI_MAX_DATA_WIDTH 1024
  `define TVIP_AXI_MAX_DATA_WIDTH 32
`endif

`endif
